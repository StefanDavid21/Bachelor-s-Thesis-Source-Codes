module audio_rom_snake (
    input wire [19:0] addr,
    output reg [7:0] data
);
    always @* begin
        case (addr)
            20'd0: data = 8'h80;
            20'd1: data = 8'h80;
            20'd2: data = 8'h80;
            20'd3: data = 8'h80;
            20'd4: data = 8'h80;
            20'd5: data = 8'h80;
            20'd6: data = 8'h80;
            20'd7: data = 8'h80;
            20'd8: data = 8'h80;
            20'd9: data = 8'h80;
            20'd10: data = 8'h80;
            20'd11: data = 8'h80;
            20'd12: data = 8'h80;
            20'd13: data = 8'h80;
            20'd14: data = 8'h80;
            20'd15: data = 8'h80;
            20'd16: data = 8'h80;
            20'd17: data = 8'h80;
            20'd18: data = 8'h80;
            20'd19: data = 8'h80;
            20'd20: data = 8'h80;
            20'd21: data = 8'h80;
            20'd22: data = 8'h80;
            20'd23: data = 8'h80;
            20'd24: data = 8'h80;
            20'd25: data = 8'h80;
            20'd26: data = 8'h80;
            20'd27: data = 8'h80;
            20'd28: data = 8'h80;
            20'd29: data = 8'h80;
            20'd30: data = 8'h80;
            20'd31: data = 8'h80;
            20'd32: data = 8'h80;
            20'd33: data = 8'h80;
            20'd34: data = 8'h80;
            20'd35: data = 8'h80;
            20'd36: data = 8'h80;
            20'd37: data = 8'h80;
            20'd38: data = 8'h80;
            20'd39: data = 8'h80;
            20'd40: data = 8'h80;
            20'd41: data = 8'h80;
            20'd42: data = 8'h80;
            20'd43: data = 8'h80;
            20'd44: data = 8'h80;
            20'd45: data = 8'h80;
            20'd46: data = 8'h80;
            20'd47: data = 8'h80;
            20'd48: data = 8'h80;
            20'd49: data = 8'h80;
            20'd50: data = 8'h80;
            20'd51: data = 8'h80;
            20'd52: data = 8'h80;
            20'd53: data = 8'h80;
            20'd54: data = 8'h80;
            20'd55: data = 8'h80;
            20'd56: data = 8'h80;
            20'd57: data = 8'h80;
            20'd58: data = 8'h80;
            20'd59: data = 8'h80;
            20'd60: data = 8'h80;
            20'd61: data = 8'h80;
            20'd62: data = 8'h80;
            20'd63: data = 8'h80;
            20'd64: data = 8'h80;
            20'd65: data = 8'h80;
            20'd66: data = 8'h80;
            20'd67: data = 8'h80;
            20'd68: data = 8'h80;
            20'd69: data = 8'h80;
            20'd70: data = 8'h80;
            20'd71: data = 8'h80;
            20'd72: data = 8'h80;
            20'd73: data = 8'h80;
            20'd74: data = 8'h80;
            20'd75: data = 8'h80;
            20'd76: data = 8'h80;
            20'd77: data = 8'h80;
            20'd78: data = 8'h80;
            20'd79: data = 8'h80;
            20'd80: data = 8'h80;
            20'd81: data = 8'h80;
            20'd82: data = 8'h80;
            20'd83: data = 8'h80;
            20'd84: data = 8'h80;
            20'd85: data = 8'h80;
            20'd86: data = 8'h80;
            20'd87: data = 8'h80;
            20'd88: data = 8'h80;
            20'd89: data = 8'h80;
            20'd90: data = 8'h80;
            20'd91: data = 8'h80;
            20'd92: data = 8'h80;
            20'd93: data = 8'h80;
            20'd94: data = 8'h80;
            20'd95: data = 8'h80;
            20'd96: data = 8'h80;
            20'd97: data = 8'h80;
            20'd98: data = 8'h80;
            20'd99: data = 8'h80;
            20'd100: data = 8'h80;
            20'd101: data = 8'h80;
            20'd102: data = 8'h80;
            20'd103: data = 8'h80;
            20'd104: data = 8'h80;
            20'd105: data = 8'h80;
            20'd106: data = 8'h80;
            20'd107: data = 8'h80;
            20'd108: data = 8'h80;
            20'd109: data = 8'h80;
            20'd110: data = 8'h80;
            20'd111: data = 8'h80;
            20'd112: data = 8'h80;
            20'd113: data = 8'h80;
            20'd114: data = 8'h80;
            20'd115: data = 8'h80;
            20'd116: data = 8'h80;
            20'd117: data = 8'h80;
            20'd118: data = 8'h80;
            20'd119: data = 8'h80;
            20'd120: data = 8'h80;
            20'd121: data = 8'h80;
            20'd122: data = 8'h80;
            20'd123: data = 8'h80;
            20'd124: data = 8'h80;
            20'd125: data = 8'h80;
            20'd126: data = 8'h80;
            20'd127: data = 8'h80;
            20'd128: data = 8'h80;
            20'd129: data = 8'h80;
            20'd130: data = 8'h80;
            20'd131: data = 8'h80;
            20'd132: data = 8'h80;
            20'd133: data = 8'h80;
            20'd134: data = 8'h80;
            20'd135: data = 8'h80;
            20'd136: data = 8'h80;
            20'd137: data = 8'h80;
            20'd138: data = 8'h80;
            20'd139: data = 8'h80;
            20'd140: data = 8'h80;
            20'd141: data = 8'h80;
            20'd142: data = 8'h80;
            20'd143: data = 8'h80;
            20'd144: data = 8'h80;
            20'd145: data = 8'h80;
            20'd146: data = 8'h80;
            20'd147: data = 8'h80;
            20'd148: data = 8'h80;
            20'd149: data = 8'h80;
            20'd150: data = 8'h80;
            20'd151: data = 8'h80;
            20'd152: data = 8'h80;
            20'd153: data = 8'h80;
            20'd154: data = 8'h80;
            20'd155: data = 8'h80;
            20'd156: data = 8'h80;
            20'd157: data = 8'h80;
            20'd158: data = 8'h80;
            20'd159: data = 8'h80;
            20'd160: data = 8'h80;
            20'd161: data = 8'h80;
            20'd162: data = 8'h80;
            20'd163: data = 8'h80;
            20'd164: data = 8'h80;
            20'd165: data = 8'h80;
            20'd166: data = 8'h80;
            20'd167: data = 8'h80;
            20'd168: data = 8'h80;
            20'd169: data = 8'h80;
            20'd170: data = 8'h80;
            20'd171: data = 8'h80;
            20'd172: data = 8'h80;
            20'd173: data = 8'h80;
            20'd174: data = 8'h80;
            20'd175: data = 8'h80;
            20'd176: data = 8'h80;
            20'd177: data = 8'h80;
            20'd178: data = 8'h80;
            20'd179: data = 8'h80;
            20'd180: data = 8'h80;
            20'd181: data = 8'h80;
            20'd182: data = 8'h80;
            20'd183: data = 8'h80;
            20'd184: data = 8'h80;
            20'd185: data = 8'h80;
            20'd186: data = 8'h80;
            20'd187: data = 8'h80;
            20'd188: data = 8'h80;
            20'd189: data = 8'h80;
            20'd190: data = 8'h80;
            20'd191: data = 8'h80;
            20'd192: data = 8'h80;
            20'd193: data = 8'h80;
            20'd194: data = 8'h80;
            20'd195: data = 8'h80;
            20'd196: data = 8'h80;
            20'd197: data = 8'h80;
            20'd198: data = 8'h80;
            20'd199: data = 8'h80;
            20'd200: data = 8'h80;
            20'd201: data = 8'h80;
            20'd202: data = 8'h80;
            20'd203: data = 8'h80;
            20'd204: data = 8'h80;
            20'd205: data = 8'h80;
            20'd206: data = 8'h80;
            20'd207: data = 8'h80;
            20'd208: data = 8'h80;
            20'd209: data = 8'h80;
            20'd210: data = 8'h80;
            20'd211: data = 8'h80;
            20'd212: data = 8'h80;
            20'd213: data = 8'h80;
            20'd214: data = 8'h80;
            20'd215: data = 8'h80;
            20'd216: data = 8'h80;
            20'd217: data = 8'h80;
            20'd218: data = 8'h80;
            20'd219: data = 8'h80;
            20'd220: data = 8'h80;
            20'd221: data = 8'h80;
            20'd222: data = 8'h80;
            20'd223: data = 8'h80;
            20'd224: data = 8'h80;
            20'd225: data = 8'h80;
            20'd226: data = 8'h80;
            20'd227: data = 8'h80;
            20'd228: data = 8'h80;
            20'd229: data = 8'h80;
            20'd230: data = 8'h80;
            20'd231: data = 8'h80;
            20'd232: data = 8'h80;
            20'd233: data = 8'h80;
            20'd234: data = 8'h80;
            20'd235: data = 8'h80;
            20'd236: data = 8'h80;
            20'd237: data = 8'h80;
            20'd238: data = 8'h80;
            20'd239: data = 8'h80;
            20'd240: data = 8'h80;
            20'd241: data = 8'h80;
            20'd242: data = 8'h80;
            20'd243: data = 8'h80;
            20'd244: data = 8'h80;
            20'd245: data = 8'h80;
            20'd246: data = 8'h80;
            20'd247: data = 8'h80;
            20'd248: data = 8'h80;
            20'd249: data = 8'h80;
            20'd250: data = 8'h80;
            20'd251: data = 8'h80;
            20'd252: data = 8'h80;
            20'd253: data = 8'h80;
            20'd254: data = 8'h80;
            20'd255: data = 8'h80;
            20'd256: data = 8'h80;
            20'd257: data = 8'h80;
            20'd258: data = 8'h80;
            20'd259: data = 8'h80;
            20'd260: data = 8'h80;
            20'd261: data = 8'h80;
            20'd262: data = 8'h80;
            20'd263: data = 8'h80;
            20'd264: data = 8'h80;
            20'd265: data = 8'h80;
            20'd266: data = 8'h80;
            20'd267: data = 8'h80;
            20'd268: data = 8'h80;
            20'd269: data = 8'h80;
            20'd270: data = 8'h80;
            20'd271: data = 8'h80;
            20'd272: data = 8'h80;
            20'd273: data = 8'h80;
            20'd274: data = 8'h80;
            20'd275: data = 8'h80;
            20'd276: data = 8'h80;
            20'd277: data = 8'h80;
            20'd278: data = 8'h80;
            20'd279: data = 8'h80;
            20'd280: data = 8'h80;
            20'd281: data = 8'h80;
            20'd282: data = 8'h80;
            20'd283: data = 8'h80;
            20'd284: data = 8'h80;
            20'd285: data = 8'h80;
            20'd286: data = 8'h80;
            20'd287: data = 8'h80;
            20'd288: data = 8'h80;
            20'd289: data = 8'h80;
            20'd290: data = 8'h80;
            20'd291: data = 8'h80;
            20'd292: data = 8'h80;
            20'd293: data = 8'h80;
            20'd294: data = 8'h80;
            20'd295: data = 8'h80;
            20'd296: data = 8'h80;
            20'd297: data = 8'h80;
            20'd298: data = 8'h80;
            20'd299: data = 8'h80;
            20'd300: data = 8'h80;
            20'd301: data = 8'h80;
            20'd302: data = 8'h80;
            20'd303: data = 8'h80;
            20'd304: data = 8'h80;
            20'd305: data = 8'h80;
            20'd306: data = 8'h80;
            20'd307: data = 8'h80;
            20'd308: data = 8'h80;
            20'd309: data = 8'h80;
            20'd310: data = 8'h80;
            20'd311: data = 8'h80;
            20'd312: data = 8'h80;
            20'd313: data = 8'h80;
            20'd314: data = 8'h80;
            20'd315: data = 8'h80;
            20'd316: data = 8'h80;
            20'd317: data = 8'h80;
            20'd318: data = 8'h80;
            20'd319: data = 8'h80;
            20'd320: data = 8'h80;
            20'd321: data = 8'h80;
            20'd322: data = 8'h80;
            20'd323: data = 8'h80;
            20'd324: data = 8'h80;
            20'd325: data = 8'h80;
            20'd326: data = 8'h80;
            20'd327: data = 8'h80;
            20'd328: data = 8'h80;
            20'd329: data = 8'h80;
            20'd330: data = 8'h80;
            20'd331: data = 8'h80;
            20'd332: data = 8'h80;
            20'd333: data = 8'h80;
            20'd334: data = 8'h80;
            20'd335: data = 8'h80;
            20'd336: data = 8'h80;
            20'd337: data = 8'h80;
            20'd338: data = 8'h80;
            20'd339: data = 8'h80;
            20'd340: data = 8'h80;
            20'd341: data = 8'h80;
            20'd342: data = 8'h80;
            20'd343: data = 8'h80;
            20'd344: data = 8'h80;
            20'd345: data = 8'h80;
            20'd346: data = 8'h80;
            20'd347: data = 8'h80;
            20'd348: data = 8'h80;
            20'd349: data = 8'h80;
            20'd350: data = 8'h80;
            20'd351: data = 8'h80;
            20'd352: data = 8'h80;
            20'd353: data = 8'h80;
            20'd354: data = 8'h80;
            20'd355: data = 8'h80;
            20'd356: data = 8'h80;
            20'd357: data = 8'h80;
            20'd358: data = 8'h80;
            20'd359: data = 8'h80;
            20'd360: data = 8'h80;
            20'd361: data = 8'h80;
            20'd362: data = 8'h80;
            20'd363: data = 8'h80;
            20'd364: data = 8'h80;
            20'd365: data = 8'h80;
            20'd366: data = 8'h80;
            20'd367: data = 8'h80;
            20'd368: data = 8'h80;
            20'd369: data = 8'h80;
            20'd370: data = 8'h80;
            20'd371: data = 8'h80;
            20'd372: data = 8'h80;
            20'd373: data = 8'h80;
            20'd374: data = 8'h80;
            20'd375: data = 8'h80;
            20'd376: data = 8'h80;
            20'd377: data = 8'h80;
            20'd378: data = 8'h80;
            20'd379: data = 8'h80;
            20'd380: data = 8'h80;
            20'd381: data = 8'h80;
            20'd382: data = 8'h80;
            20'd383: data = 8'h80;
            20'd384: data = 8'h80;
            20'd385: data = 8'h80;
            20'd386: data = 8'h80;
            20'd387: data = 8'h80;
            20'd388: data = 8'h80;
            20'd389: data = 8'h80;
            20'd390: data = 8'h80;
            20'd391: data = 8'h80;
            20'd392: data = 8'h80;
            20'd393: data = 8'h80;
            20'd394: data = 8'h80;
            20'd395: data = 8'h80;
            20'd396: data = 8'h80;
            20'd397: data = 8'h80;
            20'd398: data = 8'h80;
            20'd399: data = 8'h80;
            20'd400: data = 8'h80;
            20'd401: data = 8'h80;
            20'd402: data = 8'h80;
            20'd403: data = 8'h80;
            20'd404: data = 8'h80;
            20'd405: data = 8'h80;
            20'd406: data = 8'h80;
            20'd407: data = 8'h80;
            20'd408: data = 8'h80;
            20'd409: data = 8'h80;
            20'd410: data = 8'h80;
            20'd411: data = 8'h80;
            20'd412: data = 8'h80;
            20'd413: data = 8'h80;
            20'd414: data = 8'h80;
            20'd415: data = 8'h80;
            20'd416: data = 8'h80;
            20'd417: data = 8'h80;
            20'd418: data = 8'h80;
            20'd419: data = 8'h80;
            20'd420: data = 8'h80;
            20'd421: data = 8'h80;
            20'd422: data = 8'h80;
            20'd423: data = 8'h80;
            20'd424: data = 8'h80;
            20'd425: data = 8'h80;
            20'd426: data = 8'h7F;
            20'd427: data = 8'h7F;
            20'd428: data = 8'h80;
            20'd429: data = 8'h80;
            20'd430: data = 8'h80;
            20'd431: data = 8'h80;
            20'd432: data = 8'h80;
            20'd433: data = 8'h80;
            20'd434: data = 8'h80;
            20'd435: data = 8'h80;
            20'd436: data = 8'h80;
            20'd437: data = 8'h80;
            20'd438: data = 8'h80;
            20'd439: data = 8'h80;
            20'd440: data = 8'h80;
            20'd441: data = 8'h80;
            20'd442: data = 8'h80;
            20'd443: data = 8'h80;
            20'd444: data = 8'h80;
            20'd445: data = 8'h80;
            20'd446: data = 8'h7F;
            20'd447: data = 8'h7F;
            20'd448: data = 8'h7F;
            20'd449: data = 8'h7F;
            20'd450: data = 8'h80;
            20'd451: data = 8'h80;
            20'd452: data = 8'h7F;
            20'd453: data = 8'h7F;
            20'd454: data = 8'h80;
            20'd455: data = 8'h80;
            20'd456: data = 8'h80;
            20'd457: data = 8'h80;
            20'd458: data = 8'h7F;
            20'd459: data = 8'h7F;
            20'd460: data = 8'h80;
            20'd461: data = 8'h80;
            20'd462: data = 8'h80;
            20'd463: data = 8'h80;
            20'd464: data = 8'h80;
            20'd465: data = 8'h80;
            20'd466: data = 8'h80;
            20'd467: data = 8'h80;
            20'd468: data = 8'h7F;
            20'd469: data = 8'h7F;
            20'd470: data = 8'h80;
            20'd471: data = 8'h80;
            20'd472: data = 8'h80;
            20'd473: data = 8'h80;
            20'd474: data = 8'h7F;
            20'd475: data = 8'h7F;
            20'd476: data = 8'h80;
            20'd477: data = 8'h80;
            20'd478: data = 8'h7F;
            20'd479: data = 8'h7F;
            20'd480: data = 8'h7F;
            20'd481: data = 8'h7F;
            20'd482: data = 8'h7F;
            20'd483: data = 8'h80;
            20'd484: data = 8'h80;
            20'd485: data = 8'h80;
            20'd486: data = 8'h80;
            20'd487: data = 8'h80;
            20'd488: data = 8'h80;
            20'd489: data = 8'h80;
            20'd490: data = 8'h7F;
            20'd491: data = 8'h7F;
            20'd492: data = 8'h80;
            20'd493: data = 8'h80;
            20'd494: data = 8'h7F;
            20'd495: data = 8'h7F;
            20'd496: data = 8'h80;
            20'd497: data = 8'h80;
            20'd498: data = 8'h7F;
            20'd499: data = 8'h7F;
            20'd500: data = 8'h80;
            20'd501: data = 8'h80;
            20'd502: data = 8'h7F;
            20'd503: data = 8'h7F;
            20'd504: data = 8'h7F;
            20'd505: data = 8'h7F;
            20'd506: data = 8'h7F;
            20'd507: data = 8'h7F;
            20'd508: data = 8'h7F;
            20'd509: data = 8'h7F;
            20'd510: data = 8'h80;
            20'd511: data = 8'h80;
            20'd512: data = 8'h80;
            20'd513: data = 8'h80;
            20'd514: data = 8'h7F;
            20'd515: data = 8'h7F;
            20'd516: data = 8'h80;
            20'd517: data = 8'h80;
            20'd518: data = 8'h7F;
            20'd519: data = 8'h7F;
            20'd520: data = 8'h80;
            20'd521: data = 8'h80;
            20'd522: data = 8'h7F;
            20'd523: data = 8'h7F;
            20'd524: data = 8'h80;
            20'd525: data = 8'h80;
            20'd526: data = 8'h7F;
            20'd527: data = 8'h80;
            20'd528: data = 8'h7F;
            20'd529: data = 8'h7F;
            20'd530: data = 8'h7F;
            20'd531: data = 8'h7F;
            20'd532: data = 8'h80;
            20'd533: data = 8'h80;
            20'd534: data = 8'h80;
            20'd535: data = 8'h80;
            20'd536: data = 8'h80;
            20'd537: data = 8'h80;
            20'd538: data = 8'h7F;
            20'd539: data = 8'h7F;
            20'd540: data = 8'h80;
            20'd541: data = 8'h80;
            20'd542: data = 8'h7F;
            20'd543: data = 8'h7F;
            20'd544: data = 8'h7F;
            20'd545: data = 8'h7F;
            20'd546: data = 8'h7F;
            20'd547: data = 8'h7F;
            20'd548: data = 8'h7F;
            20'd549: data = 8'h7F;
            20'd550: data = 8'h80;
            20'd551: data = 8'h80;
            20'd552: data = 8'h80;
            20'd553: data = 8'h80;
            20'd554: data = 8'h7F;
            20'd555: data = 8'h7F;
            20'd556: data = 8'h80;
            20'd557: data = 8'h80;
            20'd558: data = 8'h7F;
            20'd559: data = 8'h7F;
            20'd560: data = 8'h80;
            20'd561: data = 8'h80;
            20'd562: data = 8'h7F;
            20'd563: data = 8'h7F;
            20'd564: data = 8'h80;
            20'd565: data = 8'h80;
            20'd566: data = 8'h7F;
            20'd567: data = 8'h7F;
            20'd568: data = 8'h80;
            20'd569: data = 8'h80;
            20'd570: data = 8'h7F;
            20'd571: data = 8'h7F;
            20'd572: data = 8'h80;
            20'd573: data = 8'h80;
            20'd574: data = 8'h7F;
            20'd575: data = 8'h7F;
            20'd576: data = 8'h80;
            20'd577: data = 8'h80;
            20'd578: data = 8'h7F;
            20'd579: data = 8'h7F;
            20'd580: data = 8'h80;
            20'd581: data = 8'h80;
            20'd582: data = 8'h7F;
            20'd583: data = 8'h7F;
            20'd584: data = 8'h80;
            20'd585: data = 8'h80;
            20'd586: data = 8'h7F;
            20'd587: data = 8'h7F;
            20'd588: data = 8'h80;
            20'd589: data = 8'h80;
            20'd590: data = 8'h80;
            20'd591: data = 8'h80;
            20'd592: data = 8'h80;
            20'd593: data = 8'h80;
            20'd594: data = 8'h80;
            20'd595: data = 8'h80;
            20'd596: data = 8'h7F;
            20'd597: data = 8'h7F;
            20'd598: data = 8'h7F;
            20'd599: data = 8'h7F;
            20'd600: data = 8'h7F;
            20'd601: data = 8'h7F;
            20'd602: data = 8'h7F;
            20'd603: data = 8'h7F;
            20'd604: data = 8'h80;
            20'd605: data = 8'h80;
            20'd606: data = 8'h7F;
            20'd607: data = 8'h7F;
            20'd608: data = 8'h7F;
            20'd609: data = 8'h7F;
            20'd610: data = 8'h80;
            20'd611: data = 8'h80;
            20'd612: data = 8'h80;
            20'd613: data = 8'h80;
            20'd614: data = 8'h80;
            20'd615: data = 8'h80;
            20'd616: data = 8'h7F;
            20'd617: data = 8'h7F;
            20'd618: data = 8'h7F;
            20'd619: data = 8'h7F;
            20'd620: data = 8'hAA;
            20'd621: data = 8'hAA;
            20'd622: data = 8'hB0;
            20'd623: data = 8'hB0;
            20'd624: data = 8'h9C;
            20'd625: data = 8'h9C;
            20'd626: data = 8'h8F;
            20'd627: data = 8'h8F;
            20'd628: data = 8'h81;
            20'd629: data = 8'h81;
            20'd630: data = 8'h79;
            20'd631: data = 8'h79;
            20'd632: data = 8'h70;
            20'd633: data = 8'h70;
            20'd634: data = 8'h6C;
            20'd635: data = 8'h6C;
            20'd636: data = 8'h69;
            20'd637: data = 8'h69;
            20'd638: data = 8'h68;
            20'd639: data = 8'h68;
            20'd640: data = 8'h6A;
            20'd641: data = 8'h6A;
            20'd642: data = 8'h6B;
            20'd643: data = 8'h6B;
            20'd644: data = 8'h6E;
            20'd645: data = 8'h6E;
            20'd646: data = 8'h59;
            20'd647: data = 8'h58;
            20'd648: data = 8'h35;
            20'd649: data = 8'h35;
            20'd650: data = 8'h4E;
            20'd651: data = 8'h4E;
            20'd652: data = 8'h63;
            20'd653: data = 8'h63;
            20'd654: data = 8'h77;
            20'd655: data = 8'h77;
            20'd656: data = 8'h85;
            20'd657: data = 8'h85;
            20'd658: data = 8'h91;
            20'd659: data = 8'h91;
            20'd660: data = 8'h99;
            20'd661: data = 8'h99;
            20'd662: data = 8'h9C;
            20'd663: data = 8'h9C;
            20'd664: data = 8'h9F;
            20'd665: data = 8'h9F;
            20'd666: data = 8'hA1;
            20'd667: data = 8'hA1;
            20'd668: data = 8'h9E;
            20'd669: data = 8'h9E;
            20'd670: data = 8'h9B;
            20'd671: data = 8'h9B;
            20'd672: data = 8'hC2;
            20'd673: data = 8'hC2;
            20'd674: data = 8'hD2;
            20'd675: data = 8'hD2;
            20'd676: data = 8'hB9;
            20'd677: data = 8'hB9;
            20'd678: data = 8'hA3;
            20'd679: data = 8'hA3;
            20'd680: data = 8'h90;
            20'd681: data = 8'h90;
            20'd682: data = 8'h7F;
            20'd683: data = 8'h7F;
            20'd684: data = 8'h73;
            20'd685: data = 8'h73;
            20'd686: data = 8'h69;
            20'd687: data = 8'h69;
            20'd688: data = 8'h64;
            20'd689: data = 8'h64;
            20'd690: data = 8'h60;
            20'd691: data = 8'h60;
            20'd692: data = 8'h5F;
            20'd693: data = 8'h5F;
            20'd694: data = 8'h60;
            20'd695: data = 8'h60;
            20'd696: data = 8'h61;
            20'd697: data = 8'h61;
            20'd698: data = 8'h29;
            20'd699: data = 8'h29;
            20'd700: data = 8'h2A;
            20'd701: data = 8'h2A;
            20'd702: data = 8'h45;
            20'd703: data = 8'h45;
            20'd704: data = 8'h5A;
            20'd705: data = 8'h5A;
            20'd706: data = 8'h6B;
            20'd707: data = 8'h6B;
            20'd708: data = 8'h7E;
            20'd709: data = 8'h7E;
            20'd710: data = 8'h8A;
            20'd711: data = 8'h8A;
            20'd712: data = 8'h94;
            20'd713: data = 8'h94;
            20'd714: data = 8'h9A;
            20'd715: data = 8'h9A;
            20'd716: data = 8'h9F;
            20'd717: data = 8'h9F;
            20'd718: data = 8'hA1;
            20'd719: data = 8'hA1;
            20'd720: data = 8'hA1;
            20'd721: data = 8'hA1;
            20'd722: data = 8'hA0;
            20'd723: data = 8'hA0;
            20'd724: data = 8'hE6;
            20'd725: data = 8'hE6;
            20'd726: data = 8'hD6;
            20'd727: data = 8'hD6;
            20'd728: data = 8'hBC;
            20'd729: data = 8'hBC;
            20'd730: data = 8'hA6;
            20'd731: data = 8'hA6;
            20'd732: data = 8'h94;
            20'd733: data = 8'h94;
            20'd734: data = 8'h84;
            20'd735: data = 8'h84;
            20'd736: data = 8'h76;
            20'd737: data = 8'h76;
            20'd738: data = 8'h6C;
            20'd739: data = 8'h6C;
            20'd740: data = 8'h67;
            20'd741: data = 8'h67;
            20'd742: data = 8'h61;
            20'd743: data = 8'h61;
            20'd744: data = 8'h5F;
            20'd745: data = 8'h5F;
            20'd746: data = 8'h5F;
            20'd747: data = 8'h5F;
            20'd748: data = 8'h5F;
            20'd749: data = 8'h5F;
            20'd750: data = 8'h10;
            20'd751: data = 8'h10;
            20'd752: data = 8'h29;
            20'd753: data = 8'h29;
            20'd754: data = 8'h45;
            20'd755: data = 8'h45;
            20'd756: data = 8'h58;
            20'd757: data = 8'h58;
            20'd758: data = 8'h6A;
            20'd759: data = 8'h6A;
            20'd760: data = 8'h7C;
            20'd761: data = 8'h7C;
            20'd762: data = 8'h87;
            20'd763: data = 8'h87;
            20'd764: data = 8'h91;
            20'd765: data = 8'h91;
            20'd766: data = 8'h97;
            20'd767: data = 8'h97;
            20'd768: data = 8'h9D;
            20'd769: data = 8'h9D;
            20'd770: data = 8'h9E;
            20'd771: data = 8'h9E;
            20'd772: data = 8'hA0;
            20'd773: data = 8'hA0;
            20'd774: data = 8'h9F;
            20'd775: data = 8'h9F;
            20'd776: data = 8'hF1;
            20'd777: data = 8'hF1;
            20'd778: data = 8'hD3;
            20'd779: data = 8'hD3;
            20'd780: data = 8'hB9;
            20'd781: data = 8'hB9;
            20'd782: data = 8'hA4;
            20'd783: data = 8'hA4;
            20'd784: data = 8'h92;
            20'd785: data = 8'h92;
            20'd786: data = 8'h82;
            20'd787: data = 8'h82;
            20'd788: data = 8'h78;
            20'd789: data = 8'h78;
            20'd790: data = 8'h6E;
            20'd791: data = 8'h6E;
            20'd792: data = 8'h68;
            20'd793: data = 8'h68;
            20'd794: data = 8'h63;
            20'd795: data = 8'h63;
            20'd796: data = 8'h62;
            20'd797: data = 8'h62;
            20'd798: data = 8'h5E;
            20'd799: data = 8'h5E;
            20'd800: data = 8'h5E;
            20'd801: data = 8'h5E;
            20'd802: data = 8'h0F;
            20'd803: data = 8'h0F;
            20'd804: data = 8'h2E;
            20'd805: data = 8'h2E;
            20'd806: data = 8'h48;
            20'd807: data = 8'h48;
            20'd808: data = 8'h5D;
            20'd809: data = 8'h5D;
            20'd810: data = 8'h6F;
            20'd811: data = 8'h6F;
            20'd812: data = 8'h7E;
            20'd813: data = 8'h7E;
            20'd814: data = 8'h89;
            20'd815: data = 8'h89;
            20'd816: data = 8'h91;
            20'd817: data = 8'h91;
            20'd818: data = 8'h97;
            20'd819: data = 8'h97;
            20'd820: data = 8'h9D;
            20'd821: data = 8'h9D;
            20'd822: data = 8'h9E;
            20'd823: data = 8'h9E;
            20'd824: data = 8'h9E;
            20'd825: data = 8'h9E;
            20'd826: data = 8'h9F;
            20'd827: data = 8'h9F;
            20'd828: data = 8'hED;
            20'd829: data = 8'hED;
            20'd830: data = 8'hCE;
            20'd831: data = 8'hCE;
            20'd832: data = 8'hB5;
            20'd833: data = 8'hB5;
            20'd834: data = 8'hA1;
            20'd835: data = 8'hA1;
            20'd836: data = 8'h8E;
            20'd837: data = 8'h8E;
            20'd838: data = 8'h81;
            20'd839: data = 8'h81;
            20'd840: data = 8'h75;
            20'd841: data = 8'h75;
            20'd842: data = 8'h6D;
            20'd843: data = 8'h6D;
            20'd844: data = 8'h67;
            20'd845: data = 8'h67;
            20'd846: data = 8'h62;
            20'd847: data = 8'h62;
            20'd848: data = 8'h61;
            20'd849: data = 8'h61;
            20'd850: data = 8'h62;
            20'd851: data = 8'h62;
            20'd852: data = 8'h63;
            20'd853: data = 8'h63;
            20'd854: data = 8'h17;
            20'd855: data = 8'h17;
            20'd856: data = 8'h35;
            20'd857: data = 8'h35;
            20'd858: data = 8'h4B;
            20'd859: data = 8'h4B;
            20'd860: data = 8'h60;
            20'd861: data = 8'h60;
            20'd862: data = 8'h72;
            20'd863: data = 8'h72;
            20'd864: data = 8'h80;
            20'd865: data = 8'h80;
            20'd866: data = 8'h8B;
            20'd867: data = 8'h8B;
            20'd868: data = 8'h93;
            20'd869: data = 8'h93;
            20'd870: data = 8'h99;
            20'd871: data = 8'h99;
            20'd872: data = 8'h9E;
            20'd873: data = 8'h9E;
            20'd874: data = 8'h9E;
            20'd875: data = 8'h9E;
            20'd876: data = 8'h9E;
            20'd877: data = 8'h9E;
            20'd878: data = 8'h9A;
            20'd879: data = 8'h9A;
            20'd880: data = 8'hE4;
            20'd881: data = 8'hE4;
            20'd882: data = 8'hC7;
            20'd883: data = 8'hC7;
            20'd884: data = 8'hB2;
            20'd885: data = 8'hB2;
            20'd886: data = 8'h9D;
            20'd887: data = 8'h9D;
            20'd888: data = 8'h8C;
            20'd889: data = 8'h8C;
            20'd890: data = 8'h7E;
            20'd891: data = 8'h7E;
            20'd892: data = 8'h73;
            20'd893: data = 8'h73;
            20'd894: data = 8'h6C;
            20'd895: data = 8'h6C;
            20'd896: data = 8'h66;
            20'd897: data = 8'h66;
            20'd898: data = 8'h62;
            20'd899: data = 8'h62;
            20'd900: data = 8'h60;
            20'd901: data = 8'h60;
            20'd902: data = 8'h60;
            20'd903: data = 8'h60;
            20'd904: data = 8'h64;
            20'd905: data = 8'h64;
            20'd906: data = 8'h1F;
            20'd907: data = 8'h1F;
            20'd908: data = 8'h39;
            20'd909: data = 8'h39;
            20'd910: data = 8'h50;
            20'd911: data = 8'h50;
            20'd912: data = 8'h63;
            20'd913: data = 8'h63;
            20'd914: data = 8'h73;
            20'd915: data = 8'h73;
            20'd916: data = 8'h82;
            20'd917: data = 8'h82;
            20'd918: data = 8'h8D;
            20'd919: data = 8'h8D;
            20'd920: data = 8'h93;
            20'd921: data = 8'h93;
            20'd922: data = 8'h99;
            20'd923: data = 8'h99;
            20'd924: data = 8'h9C;
            20'd925: data = 8'h9C;
            20'd926: data = 8'h9E;
            20'd927: data = 8'h9E;
            20'd928: data = 8'h9F;
            20'd929: data = 8'h9F;
            20'd930: data = 8'hA2;
            20'd931: data = 8'hA2;
            20'd932: data = 8'hDD;
            20'd933: data = 8'hDD;
            20'd934: data = 8'hC5;
            20'd935: data = 8'hC5;
            20'd936: data = 8'hAE;
            20'd937: data = 8'hAE;
            20'd938: data = 8'h9A;
            20'd939: data = 8'h9A;
            20'd940: data = 8'h8A;
            20'd941: data = 8'h8A;
            20'd942: data = 8'h7D;
            20'd943: data = 8'h7D;
            20'd944: data = 8'h72;
            20'd945: data = 8'h72;
            20'd946: data = 8'h6A;
            20'd947: data = 8'h6A;
            20'd948: data = 8'h66;
            20'd949: data = 8'h66;
            20'd950: data = 8'h63;
            20'd951: data = 8'h62;
            20'd952: data = 8'h60;
            20'd953: data = 8'h60;
            20'd954: data = 8'h60;
            20'd955: data = 8'h60;
            20'd956: data = 8'h52;
            20'd957: data = 8'h52;
            20'd958: data = 8'h24;
            20'd959: data = 8'h24;
            20'd960: data = 8'h3C;
            20'd961: data = 8'h3C;
            20'd962: data = 8'h53;
            20'd963: data = 8'h53;
            20'd964: data = 8'h66;
            20'd965: data = 8'h66;
            20'd966: data = 8'h75;
            20'd967: data = 8'h75;
            20'd968: data = 8'h83;
            20'd969: data = 8'h83;
            20'd970: data = 8'h8D;
            20'd971: data = 8'h8D;
            20'd972: data = 8'h95;
            20'd973: data = 8'h95;
            20'd974: data = 8'h9A;
            20'd975: data = 8'h9A;
            20'd976: data = 8'h9D;
            20'd977: data = 8'h9D;
            20'd978: data = 8'h9E;
            20'd979: data = 8'h9E;
            20'd980: data = 8'h9E;
            20'd981: data = 8'h9E;
            20'd982: data = 8'hBC;
            20'd983: data = 8'hBC;
            20'd984: data = 8'hD8;
            20'd985: data = 8'hD8;
            20'd986: data = 8'hC0;
            20'd987: data = 8'hC0;
            20'd988: data = 8'hAB;
            20'd989: data = 8'hAB;
            20'd990: data = 8'h96;
            20'd991: data = 8'h96;
            20'd992: data = 8'h87;
            20'd993: data = 8'h87;
            20'd994: data = 8'h7B;
            20'd995: data = 8'h7B;
            20'd996: data = 8'h72;
            20'd997: data = 8'h72;
            20'd998: data = 8'h6A;
            20'd999: data = 8'h6A;
            20'd1000: data = 8'h64;
            20'd1001: data = 8'h64;
            20'd1002: data = 8'h62;
            20'd1003: data = 8'h62;
            20'd1004: data = 8'h62;
            20'd1005: data = 8'h62;
            20'd1006: data = 8'h61;
            20'd1007: data = 8'h61;
            20'd1008: data = 8'h30;
            20'd1009: data = 8'h30;
            20'd1010: data = 8'h28;
            20'd1011: data = 8'h28;
            20'd1012: data = 8'h40;
            20'd1013: data = 8'h40;
            20'd1014: data = 8'h56;
            20'd1015: data = 8'h56;
            20'd1016: data = 8'h69;
            20'd1017: data = 8'h69;
            20'd1018: data = 8'h79;
            20'd1019: data = 8'h79;
            20'd1020: data = 8'h85;
            20'd1021: data = 8'h85;
            20'd1022: data = 8'h8F;
            20'd1023: data = 8'h8F;
            20'd1024: data = 8'h96;
            20'd1025: data = 8'h96;
            20'd1026: data = 8'h9A;
            20'd1027: data = 8'h9A;
            20'd1028: data = 8'h9D;
            20'd1029: data = 8'h9D;
            20'd1030: data = 8'h9E;
            20'd1031: data = 8'h9E;
            20'd1032: data = 8'h9E;
            20'd1033: data = 8'h9E;
            20'd1034: data = 8'hDF;
            20'd1035: data = 8'hDF;
            20'd1036: data = 8'hD6;
            20'd1037: data = 8'hD5;
            20'd1038: data = 8'hBD;
            20'd1039: data = 8'hBD;
            20'd1040: data = 8'hA8;
            20'd1041: data = 8'hA8;
            20'd1042: data = 8'h94;
            20'd1043: data = 8'h94;
            20'd1044: data = 8'h86;
            20'd1045: data = 8'h86;
            20'd1046: data = 8'h79;
            20'd1047: data = 8'h79;
            20'd1048: data = 8'h6F;
            20'd1049: data = 8'h6F;
            20'd1050: data = 8'h69;
            20'd1051: data = 8'h69;
            20'd1052: data = 8'h65;
            20'd1053: data = 8'h65;
            20'd1054: data = 8'h62;
            20'd1055: data = 8'h62;
            20'd1056: data = 8'h61;
            20'd1057: data = 8'h61;
            20'd1058: data = 8'h60;
            20'd1059: data = 8'h60;
            20'd1060: data = 8'h14;
            20'd1061: data = 8'h14;
            20'd1062: data = 8'h2B;
            20'd1063: data = 8'h2B;
            20'd1064: data = 8'h45;
            20'd1065: data = 8'h44;
            20'd1066: data = 8'h59;
            20'd1067: data = 8'h59;
            20'd1068: data = 8'h6C;
            20'd1069: data = 8'h6C;
            20'd1070: data = 8'h7A;
            20'd1071: data = 8'h7A;
            20'd1072: data = 8'h87;
            20'd1073: data = 8'h87;
            20'd1074: data = 8'h90;
            20'd1075: data = 8'h90;
            20'd1076: data = 8'h96;
            20'd1077: data = 8'h96;
            20'd1078: data = 8'h9B;
            20'd1079: data = 8'h9B;
            20'd1080: data = 8'h9E;
            20'd1081: data = 8'h9E;
            20'd1082: data = 8'h9E;
            20'd1083: data = 8'h9E;
            20'd1084: data = 8'h9F;
            20'd1085: data = 8'h9F;
            20'd1086: data = 8'hF1;
            20'd1087: data = 8'hF1;
            20'd1088: data = 8'hD2;
            20'd1089: data = 8'hD2;
            20'd1090: data = 8'hB8;
            20'd1091: data = 8'hB8;
            20'd1092: data = 8'hA3;
            20'd1093: data = 8'hA3;
            20'd1094: data = 8'h92;
            20'd1095: data = 8'h92;
            20'd1096: data = 8'h84;
            20'd1097: data = 8'h84;
            20'd1098: data = 8'h77;
            20'd1099: data = 8'h77;
            20'd1100: data = 8'h6E;
            20'd1101: data = 8'h6E;
            20'd1102: data = 8'h67;
            20'd1103: data = 8'h67;
            20'd1104: data = 8'h63;
            20'd1105: data = 8'h63;
            20'd1106: data = 8'h62;
            20'd1107: data = 8'h62;
            20'd1108: data = 8'h61;
            20'd1109: data = 8'h61;
            20'd1110: data = 8'h5F;
            20'd1111: data = 8'h5F;
            20'd1112: data = 8'h0E;
            20'd1113: data = 8'h0E;
            20'd1114: data = 8'h2F;
            20'd1115: data = 8'h2F;
            20'd1116: data = 8'h48;
            20'd1117: data = 8'h48;
            20'd1118: data = 8'h5D;
            20'd1119: data = 8'h5E;
            20'd1120: data = 8'h6D;
            20'd1121: data = 8'h6D;
            20'd1122: data = 8'h7E;
            20'd1123: data = 8'h7E;
            20'd1124: data = 8'h89;
            20'd1125: data = 8'h89;
            20'd1126: data = 8'h91;
            20'd1127: data = 8'h91;
            20'd1128: data = 8'h97;
            20'd1129: data = 8'h97;
            20'd1130: data = 8'h9B;
            20'd1131: data = 8'h9B;
            20'd1132: data = 8'h9D;
            20'd1133: data = 8'h9E;
            20'd1134: data = 8'h9E;
            20'd1135: data = 8'h9E;
            20'd1136: data = 8'hA0;
            20'd1137: data = 8'hA0;
            20'd1138: data = 8'hEE;
            20'd1139: data = 8'hEE;
            20'd1140: data = 8'hCE;
            20'd1141: data = 8'hCE;
            20'd1142: data = 8'hB7;
            20'd1143: data = 8'hB7;
            20'd1144: data = 8'hA0;
            20'd1145: data = 8'hA0;
            20'd1146: data = 8'h8F;
            20'd1147: data = 8'h8F;
            20'd1148: data = 8'h80;
            20'd1149: data = 8'h80;
            20'd1150: data = 8'h77;
            20'd1151: data = 8'h77;
            20'd1152: data = 8'h6E;
            20'd1153: data = 8'h6E;
            20'd1154: data = 8'h66;
            20'd1155: data = 8'h66;
            20'd1156: data = 8'h63;
            20'd1157: data = 8'h63;
            20'd1158: data = 8'h63;
            20'd1159: data = 8'h63;
            20'd1160: data = 8'h61;
            20'd1161: data = 8'h61;
            20'd1162: data = 8'h60;
            20'd1163: data = 8'h60;
            20'd1164: data = 8'h15;
            20'd1165: data = 8'h15;
            20'd1166: data = 8'h34;
            20'd1167: data = 8'h34;
            20'd1168: data = 8'h4A;
            20'd1169: data = 8'h4A;
            20'd1170: data = 8'h60;
            20'd1171: data = 8'h60;
            20'd1172: data = 8'h70;
            20'd1173: data = 8'h70;
            20'd1174: data = 8'h7F;
            20'd1175: data = 8'h7F;
            20'd1176: data = 8'h89;
            20'd1177: data = 8'h89;
            20'd1178: data = 8'h92;
            20'd1179: data = 8'h92;
            20'd1180: data = 8'h98;
            20'd1181: data = 8'h98;
            20'd1182: data = 8'h9C;
            20'd1183: data = 8'h9C;
            20'd1184: data = 8'h9D;
            20'd1185: data = 8'h9D;
            20'd1186: data = 8'h9D;
            20'd1187: data = 8'h9D;
            20'd1188: data = 8'h9C;
            20'd1189: data = 8'h9C;
            20'd1190: data = 8'hE6;
            20'd1191: data = 8'hE6;
            20'd1192: data = 8'hC8;
            20'd1193: data = 8'hC8;
            20'd1194: data = 8'hB3;
            20'd1195: data = 8'hB3;
            20'd1196: data = 8'h9E;
            20'd1197: data = 8'h9E;
            20'd1198: data = 8'h8F;
            20'd1199: data = 8'h8F;
            20'd1200: data = 8'h7F;
            20'd1201: data = 8'h7F;
            20'd1202: data = 8'h75;
            20'd1203: data = 8'h75;
            20'd1204: data = 8'h6D;
            20'd1205: data = 8'h6D;
            20'd1206: data = 8'h67;
            20'd1207: data = 8'h67;
            20'd1208: data = 8'h63;
            20'd1209: data = 8'h63;
            20'd1210: data = 8'h61;
            20'd1211: data = 8'h61;
            20'd1212: data = 8'h61;
            20'd1213: data = 8'h61;
            20'd1214: data = 8'h64;
            20'd1215: data = 8'h64;
            20'd1216: data = 8'h1D;
            20'd1217: data = 8'h1D;
            20'd1218: data = 8'h38;
            20'd1219: data = 8'h38;
            20'd1220: data = 8'h4D;
            20'd1221: data = 8'h4D;
            20'd1222: data = 8'h62;
            20'd1223: data = 8'h62;
            20'd1224: data = 8'h72;
            20'd1225: data = 8'h72;
            20'd1226: data = 8'h81;
            20'd1227: data = 8'h81;
            20'd1228: data = 8'h8C;
            20'd1229: data = 8'h8C;
            20'd1230: data = 8'h94;
            20'd1231: data = 8'h94;
            20'd1232: data = 8'h99;
            20'd1233: data = 8'h99;
            20'd1234: data = 8'h9C;
            20'd1235: data = 8'h9C;
            20'd1236: data = 8'h9F;
            20'd1237: data = 8'h9F;
            20'd1238: data = 8'h9F;
            20'd1239: data = 8'h9F;
            20'd1240: data = 8'h9D;
            20'd1241: data = 8'h9D;
            20'd1242: data = 8'hE0;
            20'd1243: data = 8'hE0;
            20'd1244: data = 8'hC6;
            20'd1245: data = 8'hC6;
            20'd1246: data = 8'hAF;
            20'd1247: data = 8'hAF;
            20'd1248: data = 8'h9A;
            20'd1249: data = 8'h9A;
            20'd1250: data = 8'h8C;
            20'd1251: data = 8'h8C;
            20'd1252: data = 8'h7E;
            20'd1253: data = 8'h7E;
            20'd1254: data = 8'h72;
            20'd1255: data = 8'h72;
            20'd1256: data = 8'h6B;
            20'd1257: data = 8'h6B;
            20'd1258: data = 8'h65;
            20'd1259: data = 8'h65;
            20'd1260: data = 8'h64;
            20'd1261: data = 8'h64;
            20'd1262: data = 8'h60;
            20'd1263: data = 8'h60;
            20'd1264: data = 8'h60;
            20'd1265: data = 8'h60;
            20'd1266: data = 8'h5A;
            20'd1267: data = 8'h5A;
            20'd1268: data = 8'h22;
            20'd1269: data = 8'h22;
            20'd1270: data = 8'h3A;
            20'd1271: data = 8'h3A;
            20'd1272: data = 8'h51;
            20'd1273: data = 8'h51;
            20'd1274: data = 8'h66;
            20'd1275: data = 8'h66;
            20'd1276: data = 8'h76;
            20'd1277: data = 8'h76;
            20'd1278: data = 8'h82;
            20'd1279: data = 8'h82;
            20'd1280: data = 8'h8D;
            20'd1281: data = 8'h8D;
            20'd1282: data = 8'h95;
            20'd1283: data = 8'h95;
            20'd1284: data = 8'h9B;
            20'd1285: data = 8'h9B;
            20'd1286: data = 8'h9C;
            20'd1287: data = 8'h9C;
            20'd1288: data = 8'h9D;
            20'd1289: data = 8'h9D;
            20'd1290: data = 8'h9F;
            20'd1291: data = 8'h9F;
            20'd1292: data = 8'hB3;
            20'd1293: data = 8'hB3;
            20'd1294: data = 8'hDA;
            20'd1295: data = 8'hDA;
            20'd1296: data = 8'hC2;
            20'd1297: data = 8'hC2;
            20'd1298: data = 8'hAB;
            20'd1299: data = 8'hAB;
            20'd1300: data = 8'h98;
            20'd1301: data = 8'h98;
            20'd1302: data = 8'h88;
            20'd1303: data = 8'h88;
            20'd1304: data = 8'h7B;
            20'd1305: data = 8'h7B;
            20'd1306: data = 8'h71;
            20'd1307: data = 8'h71;
            20'd1308: data = 8'h69;
            20'd1309: data = 8'h69;
            20'd1310: data = 8'h64;
            20'd1311: data = 8'h64;
            20'd1312: data = 8'h62;
            20'd1313: data = 8'h62;
            20'd1314: data = 8'h62;
            20'd1315: data = 8'h62;
            20'd1316: data = 8'h62;
            20'd1317: data = 8'h62;
            20'd1318: data = 8'h3A;
            20'd1319: data = 8'h3A;
            20'd1320: data = 8'h28;
            20'd1321: data = 8'h28;
            20'd1322: data = 8'h3F;
            20'd1323: data = 8'h3F;
            20'd1324: data = 8'h55;
            20'd1325: data = 8'h55;
            20'd1326: data = 8'h68;
            20'd1327: data = 8'h68;
            20'd1328: data = 8'h78;
            20'd1329: data = 8'h78;
            20'd1330: data = 8'h85;
            20'd1331: data = 8'h85;
            20'd1332: data = 8'h8E;
            20'd1333: data = 8'h8E;
            20'd1334: data = 8'h96;
            20'd1335: data = 8'h96;
            20'd1336: data = 8'h9B;
            20'd1337: data = 8'h9B;
            20'd1338: data = 8'h9D;
            20'd1339: data = 8'h9D;
            20'd1340: data = 8'h9E;
            20'd1341: data = 8'h9E;
            20'd1342: data = 8'h9D;
            20'd1343: data = 8'h9D;
            20'd1344: data = 8'hD8;
            20'd1345: data = 8'hD8;
            20'd1346: data = 8'hD6;
            20'd1347: data = 8'hD6;
            20'd1348: data = 8'hBD;
            20'd1349: data = 8'hBD;
            20'd1350: data = 8'h67;
            20'd1351: data = 8'h67;
            20'd1352: data = 8'h6D;
            20'd1353: data = 8'h6D;
            20'd1354: data = 8'h6E;
            20'd1355: data = 8'h6E;
            20'd1356: data = 8'h6F;
            20'd1357: data = 8'h6F;
            20'd1358: data = 8'h72;
            20'd1359: data = 8'h72;
            20'd1360: data = 8'h73;
            20'd1361: data = 8'h74;
            20'd1362: data = 8'h75;
            20'd1363: data = 8'h75;
            20'd1364: data = 8'h76;
            20'd1365: data = 8'h76;
            20'd1366: data = 8'h77;
            20'd1367: data = 8'h77;
            20'd1368: data = 8'h77;
            20'd1369: data = 8'h77;
            20'd1370: data = 8'h77;
            20'd1371: data = 8'h77;
            20'd1372: data = 8'h77;
            20'd1373: data = 8'h77;
            20'd1374: data = 8'h77;
            20'd1375: data = 8'h77;
            20'd1376: data = 8'h77;
            20'd1377: data = 8'h77;
            20'd1378: data = 8'h77;
            20'd1379: data = 8'h77;
            20'd1380: data = 8'h77;
            20'd1381: data = 8'h77;
            20'd1382: data = 8'h79;
            20'd1383: data = 8'h79;
            20'd1384: data = 8'h7A;
            20'd1385: data = 8'h7A;
            20'd1386: data = 8'h7C;
            20'd1387: data = 8'h7C;
            20'd1388: data = 8'h7E;
            20'd1389: data = 8'h7E;
            20'd1390: data = 8'h80;
            20'd1391: data = 8'h80;
            20'd1392: data = 8'h82;
            20'd1393: data = 8'h82;
            20'd1394: data = 8'h84;
            20'd1395: data = 8'h84;
            20'd1396: data = 8'h86;
            20'd1397: data = 8'h86;
            20'd1398: data = 8'h87;
            20'd1399: data = 8'h87;
            20'd1400: data = 8'h87;
            20'd1401: data = 8'h87;
            20'd1402: data = 8'h88;
            20'd1403: data = 8'h88;
            20'd1404: data = 8'h87;
            20'd1405: data = 8'h87;
            20'd1406: data = 8'h86;
            20'd1407: data = 8'h86;
            20'd1408: data = 8'h85;
            20'd1409: data = 8'h85;
            20'd1410: data = 8'h84;
            20'd1411: data = 8'h84;
            20'd1412: data = 8'h82;
            20'd1413: data = 8'h82;
            20'd1414: data = 8'h81;
            20'd1415: data = 8'h81;
            20'd1416: data = 8'h7F;
            20'd1417: data = 8'h7F;
            20'd1418: data = 8'h7E;
            20'd1419: data = 8'h7E;
            20'd1420: data = 8'h7D;
            20'd1421: data = 8'h7D;
            20'd1422: data = 8'h7D;
            20'd1423: data = 8'h7D;
            20'd1424: data = 8'h7C;
            20'd1425: data = 8'h7C;
            20'd1426: data = 8'h7C;
            20'd1427: data = 8'h7C;
            20'd1428: data = 8'h7C;
            20'd1429: data = 8'h7C;
            20'd1430: data = 8'h7C;
            20'd1431: data = 8'h7C;
            20'd1432: data = 8'h7D;
            20'd1433: data = 8'h7D;
            20'd1434: data = 8'h7D;
            20'd1435: data = 8'h7D;
            20'd1436: data = 8'h7D;
            20'd1437: data = 8'h7D;
            20'd1438: data = 8'h7E;
            20'd1439: data = 8'h7E;
            20'd1440: data = 8'h7E;
            20'd1441: data = 8'h7E;
            20'd1442: data = 8'h7E;
            20'd1443: data = 8'h7E;
            20'd1444: data = 8'h7E;
            20'd1445: data = 8'h7E;
            20'd1446: data = 8'h7F;
            20'd1447: data = 8'h7F;
            20'd1448: data = 8'h7F;
            20'd1449: data = 8'h7F;
            20'd1450: data = 8'h7F;
            20'd1451: data = 8'h7F;
            20'd1452: data = 8'h80;
            20'd1453: data = 8'h80;
            20'd1454: data = 8'h80;
            20'd1455: data = 8'h80;
            20'd1456: data = 8'h80;
            20'd1457: data = 8'h80;
            20'd1458: data = 8'h80;
            20'd1459: data = 8'h80;
            20'd1460: data = 8'h81;
            20'd1461: data = 8'h81;
            20'd1462: data = 8'h81;
            20'd1463: data = 8'h81;
            20'd1464: data = 8'h81;
            20'd1465: data = 8'h81;
            20'd1466: data = 8'h81;
            20'd1467: data = 8'h81;
            20'd1468: data = 8'h81;
            20'd1469: data = 8'h81;
            20'd1470: data = 8'h81;
            20'd1471: data = 8'h81;
            20'd1472: data = 8'h81;
            20'd1473: data = 8'h81;
            20'd1474: data = 8'h80;
            20'd1475: data = 8'h80;
            20'd1476: data = 8'h80;
            20'd1477: data = 8'h80;
            20'd1478: data = 8'h80;
            20'd1479: data = 8'h80;
            20'd1480: data = 8'h80;
            20'd1481: data = 8'h80;
            20'd1482: data = 8'h7F;
            20'd1483: data = 8'h7F;
            20'd1484: data = 8'h7F;
            20'd1485: data = 8'h7F;
            20'd1486: data = 8'h7F;
            20'd1487: data = 8'h7F;
            20'd1488: data = 8'h7F;
            20'd1489: data = 8'h7F;
            20'd1490: data = 8'h7F;
            20'd1491: data = 8'h7F;
            20'd1492: data = 8'h7F;
            20'd1493: data = 8'h7F;
            20'd1494: data = 8'h7F;
            20'd1495: data = 8'h7F;
            20'd1496: data = 8'h7F;
            20'd1497: data = 8'h7F;
            20'd1498: data = 8'h7F;
            20'd1499: data = 8'h7F;
            20'd1500: data = 8'h7F;
            20'd1501: data = 8'h7F;
            20'd1502: data = 8'h7F;
            20'd1503: data = 8'h7F;
            20'd1504: data = 8'h7F;
            20'd1505: data = 8'h7F;
            20'd1506: data = 8'h7F;
            20'd1507: data = 8'h7F;
            20'd1508: data = 8'h7F;
            20'd1509: data = 8'h7F;
            20'd1510: data = 8'h7F;
            20'd1511: data = 8'h7F;
            20'd1512: data = 8'h7F;
            20'd1513: data = 8'h7F;
            20'd1514: data = 8'h7F;
            20'd1515: data = 8'h7F;
            20'd1516: data = 8'h7F;
            20'd1517: data = 8'h7F;
            20'd1518: data = 8'h80;
            20'd1519: data = 8'h80;
            20'd1520: data = 8'h80;
            20'd1521: data = 8'h80;
            20'd1522: data = 8'h80;
            20'd1523: data = 8'h80;
            20'd1524: data = 8'h80;
            20'd1525: data = 8'h80;
            20'd1526: data = 8'h80;
            20'd1527: data = 8'h80;
            20'd1528: data = 8'h80;
            20'd1529: data = 8'h80;
            20'd1530: data = 8'h80;
            20'd1531: data = 8'h80;
            20'd1532: data = 8'h80;
            20'd1533: data = 8'h80;
            20'd1534: data = 8'h80;
            20'd1535: data = 8'h80;
            20'd1536: data = 8'h80;
            20'd1537: data = 8'h80;
            20'd1538: data = 8'h80;
            20'd1539: data = 8'h80;
            20'd1540: data = 8'h80;
            20'd1541: data = 8'h80;
            20'd1542: data = 8'h80;
            20'd1543: data = 8'h80;
            20'd1544: data = 8'h80;
            20'd1545: data = 8'h80;
            20'd1546: data = 8'h7F;
            20'd1547: data = 8'h7F;
            20'd1548: data = 8'h7F;
            20'd1549: data = 8'h7F;
            20'd1550: data = 8'h7F;
            20'd1551: data = 8'h7F;
            20'd1552: data = 8'h7F;
            20'd1553: data = 8'h7F;
            20'd1554: data = 8'h7F;
            20'd1555: data = 8'h7F;
            20'd1556: data = 8'h7F;
            20'd1557: data = 8'h7F;
            20'd1558: data = 8'h7F;
            20'd1559: data = 8'h7F;
            20'd1560: data = 8'h7F;
            20'd1561: data = 8'h7F;
            20'd1562: data = 8'h7F;
            20'd1563: data = 8'h7F;
            20'd1564: data = 8'h7F;
            20'd1565: data = 8'h7F;
            20'd1566: data = 8'h7F;
            20'd1567: data = 8'h7F;
            20'd1568: data = 8'h7F;
            20'd1569: data = 8'h7F;
            20'd1570: data = 8'h7F;
            20'd1571: data = 8'h7F;
            20'd1572: data = 8'h7F;
            20'd1573: data = 8'h7F;
            20'd1574: data = 8'h7F;
            20'd1575: data = 8'h7F;
            20'd1576: data = 8'h7F;
            20'd1577: data = 8'h80;
            20'd1578: data = 8'h80;
            20'd1579: data = 8'h80;
            20'd1580: data = 8'h80;
            20'd1581: data = 8'h80;
            20'd1582: data = 8'h80;
            20'd1583: data = 8'h80;
            20'd1584: data = 8'h80;
            20'd1585: data = 8'h80;
            20'd1586: data = 8'h80;
            20'd1587: data = 8'h80;
            20'd1588: data = 8'h80;
            20'd1589: data = 8'h80;
            20'd1590: data = 8'h80;
            20'd1591: data = 8'h80;
            20'd1592: data = 8'h80;
            20'd1593: data = 8'h80;
            20'd1594: data = 8'h80;
            20'd1595: data = 8'h80;
            20'd1596: data = 8'h80;
            20'd1597: data = 8'h80;
            20'd1598: data = 8'h80;
            20'd1599: data = 8'h80;
            20'd1600: data = 8'h80;
            20'd1601: data = 8'h80;
            20'd1602: data = 8'h80;
            20'd1603: data = 8'h80;
            20'd1604: data = 8'h80;
            20'd1605: data = 8'h80;
            20'd1606: data = 8'h7F;
            20'd1607: data = 8'h7F;
            20'd1608: data = 8'h7F;
            20'd1609: data = 8'h7F;
            20'd1610: data = 8'h80;
            20'd1611: data = 8'h80;
            20'd1612: data = 8'h7F;
            20'd1613: data = 8'h80;
            20'd1614: data = 8'h7F;
            20'd1615: data = 8'h80;
            20'd1616: data = 8'h80;
            20'd1617: data = 8'h7F;
            20'd1618: data = 8'h7F;
            20'd1619: data = 8'h7F;
            20'd1620: data = 8'h80;
            20'd1621: data = 8'h7F;
            20'd1622: data = 8'h80;
            20'd1623: data = 8'h7F;
            20'd1624: data = 8'h7F;
            20'd1625: data = 8'h7F;
            20'd1626: data = 8'h80;
            20'd1627: data = 8'h7F;
            20'd1628: data = 8'h7F;
            20'd1629: data = 8'h80;
            20'd1630: data = 8'h7F;
            20'd1631: data = 8'h7F;
            20'd1632: data = 8'h7F;
            20'd1633: data = 8'h80;
            20'd1634: data = 8'h7F;
            20'd1635: data = 8'h7F;
            20'd1636: data = 8'h80;
            20'd1637: data = 8'h80;
            20'd1638: data = 8'h80;
            20'd1639: data = 8'h80;
            20'd1640: data = 8'h80;
            20'd1641: data = 8'h80;
            20'd1642: data = 8'h80;
            20'd1643: data = 8'h80;
            20'd1644: data = 8'h80;
            20'd1645: data = 8'h80;
            20'd1646: data = 8'h7F;
            20'd1647: data = 8'h80;
            20'd1648: data = 8'h80;
            20'd1649: data = 8'h80;
            20'd1650: data = 8'h80;
            20'd1651: data = 8'h7F;
            20'd1652: data = 8'h80;
            20'd1653: data = 8'h80;
            20'd1654: data = 8'h80;
            20'd1655: data = 8'h80;
            20'd1656: data = 8'h80;
            20'd1657: data = 8'h80;
            20'd1658: data = 8'h80;
            20'd1659: data = 8'h80;
            20'd1660: data = 8'h80;
            20'd1661: data = 8'h80;
            20'd1662: data = 8'h80;
            20'd1663: data = 8'h80;
            20'd1664: data = 8'h7F;
            20'd1665: data = 8'h80;
            20'd1666: data = 8'h7F;
            20'd1667: data = 8'h7F;
            20'd1668: data = 8'h7F;
            20'd1669: data = 8'h80;
            20'd1670: data = 8'h7F;
            20'd1671: data = 8'h7F;
            20'd1672: data = 8'h80;
            20'd1673: data = 8'h80;
            20'd1674: data = 8'h7F;
            20'd1675: data = 8'h80;
            20'd1676: data = 8'h80;
            20'd1677: data = 8'h80;
            20'd1678: data = 8'h7F;
            20'd1679: data = 8'h7F;
            20'd1680: data = 8'h7F;
            20'd1681: data = 8'h7F;
            20'd1682: data = 8'h80;
            20'd1683: data = 8'h80;
            20'd1684: data = 8'h80;
            20'd1685: data = 8'h7F;
            20'd1686: data = 8'h80;
            20'd1687: data = 8'h80;
            20'd1688: data = 8'h80;
            20'd1689: data = 8'h7F;
            20'd1690: data = 8'h80;
            20'd1691: data = 8'h80;
            20'd1692: data = 8'h7F;
            20'd1693: data = 8'h80;
            20'd1694: data = 8'h80;
            20'd1695: data = 8'h80;
            20'd1696: data = 8'h80;
            20'd1697: data = 8'h7F;
            20'd1698: data = 8'h7F;
            20'd1699: data = 8'h80;
            20'd1700: data = 8'h80;
            20'd1701: data = 8'h80;
            20'd1702: data = 8'h80;
            20'd1703: data = 8'h80;
            20'd1704: data = 8'h7F;
            20'd1705: data = 8'h80;
            20'd1706: data = 8'h7F;
            20'd1707: data = 8'h80;
            20'd1708: data = 8'h80;
            20'd1709: data = 8'h80;
            20'd1710: data = 8'h80;
            20'd1711: data = 8'h80;
            20'd1712: data = 8'h80;
            20'd1713: data = 8'h80;
            20'd1714: data = 8'h80;
            20'd1715: data = 8'h80;
            20'd1716: data = 8'h80;
            20'd1717: data = 8'h80;
            20'd1718: data = 8'h80;
            20'd1719: data = 8'h80;
            20'd1720: data = 8'h80;
            20'd1721: data = 8'h80;
            20'd1722: data = 8'h80;
            20'd1723: data = 8'h80;
            20'd1724: data = 8'h7F;
            20'd1725: data = 8'h7F;
            20'd1726: data = 8'h80;
            20'd1727: data = 8'h80;
            20'd1728: data = 8'h80;
            20'd1729: data = 8'h80;
            20'd1730: data = 8'h80;
            20'd1731: data = 8'h80;
            20'd1732: data = 8'h7F;
            20'd1733: data = 8'h80;
            20'd1734: data = 8'h7F;
            20'd1735: data = 8'h7F;
            20'd1736: data = 8'h7F;
            20'd1737: data = 8'h80;
            20'd1738: data = 8'h80;
            20'd1739: data = 8'h80;
            20'd1740: data = 8'h80;
            20'd1741: data = 8'h80;
            20'd1742: data = 8'h7F;
            20'd1743: data = 8'h7F;
            20'd1744: data = 8'h80;
            20'd1745: data = 8'h80;
            20'd1746: data = 8'h80;
            20'd1747: data = 8'h7F;
            20'd1748: data = 8'h80;
            20'd1749: data = 8'h80;
            20'd1750: data = 8'h7F;
            20'd1751: data = 8'h80;
            20'd1752: data = 8'h80;
            20'd1753: data = 8'h80;
            20'd1754: data = 8'h7F;
            20'd1755: data = 8'h7F;
            20'd1756: data = 8'h7F;
            20'd1757: data = 8'h7F;
            20'd1758: data = 8'h80;
            20'd1759: data = 8'h80;
            20'd1760: data = 8'h80;
            20'd1761: data = 8'h7F;
            20'd1762: data = 8'h80;
            20'd1763: data = 8'h7F;
            20'd1764: data = 8'h7F;
            20'd1765: data = 8'h7F;
            20'd1766: data = 8'h7F;
            20'd1767: data = 8'h7F;
            20'd1768: data = 8'h80;
            20'd1769: data = 8'h80;
            20'd1770: data = 8'h80;
            20'd1771: data = 8'h80;
            20'd1772: data = 8'h7F;
            20'd1773: data = 8'h7F;
            20'd1774: data = 8'h7F;
            20'd1775: data = 8'h7F;
            20'd1776: data = 8'h80;
            20'd1777: data = 8'h80;
            20'd1778: data = 8'h80;
            20'd1779: data = 8'h80;
            20'd1780: data = 8'h7F;
            20'd1781: data = 8'h7F;
            20'd1782: data = 8'h7F;
            20'd1783: data = 8'h7F;
            20'd1784: data = 8'h80;
            20'd1785: data = 8'h80;
            20'd1786: data = 8'h7F;
            20'd1787: data = 8'h7F;
            20'd1788: data = 8'h80;
            20'd1789: data = 8'h80;
            20'd1790: data = 8'h7F;
            20'd1791: data = 8'h7F;
            20'd1792: data = 8'h80;
            20'd1793: data = 8'h80;
            20'd1794: data = 8'h7F;
            20'd1795: data = 8'h7F;
            20'd1796: data = 8'h80;
            20'd1797: data = 8'h80;
            20'd1798: data = 8'h7F;
            20'd1799: data = 8'h7F;
            20'd1800: data = 8'h7F;
            20'd1801: data = 8'h7F;
            20'd1802: data = 8'h80;
            20'd1803: data = 8'h80;
            20'd1804: data = 8'h80;
            20'd1805: data = 8'h80;
            20'd1806: data = 8'h7F;
            20'd1807: data = 8'h7F;
            20'd1808: data = 8'h7F;
            20'd1809: data = 8'h7F;
            20'd1810: data = 8'h7F;
            20'd1811: data = 8'h7F;
            20'd1812: data = 8'h7F;
            20'd1813: data = 8'h7F;
            20'd1814: data = 8'h80;
            20'd1815: data = 8'h80;
            20'd1816: data = 8'h7F;
            20'd1817: data = 8'h7F;
            20'd1818: data = 8'h80;
            20'd1819: data = 8'h80;
            20'd1820: data = 8'h7F;
            20'd1821: data = 8'h7F;
            20'd1822: data = 8'h80;
            20'd1823: data = 8'h80;
            20'd1824: data = 8'h80;
            20'd1825: data = 8'h80;
            20'd1826: data = 8'h80;
            20'd1827: data = 8'h7F;
            20'd1828: data = 8'h80;
            20'd1829: data = 8'h80;
            20'd1830: data = 8'h80;
            20'd1831: data = 8'h80;
            20'd1832: data = 8'h7F;
            20'd1833: data = 8'h7F;
            20'd1834: data = 8'h80;
            20'd1835: data = 8'h80;
            20'd1836: data = 8'h80;
            20'd1837: data = 8'h80;
            20'd1838: data = 8'h80;
            20'd1839: data = 8'h80;
            20'd1840: data = 8'h7F;
            20'd1841: data = 8'h80;
            20'd1842: data = 8'h7F;
            20'd1843: data = 8'h7F;
            20'd1844: data = 8'h80;
            20'd1845: data = 8'h80;
            20'd1846: data = 8'h7F;
            20'd1847: data = 8'h7F;
            20'd1848: data = 8'h7F;
            20'd1849: data = 8'h7F;
            20'd1850: data = 8'h80;
            20'd1851: data = 8'h80;
            20'd1852: data = 8'h80;
            20'd1853: data = 8'h80;
            20'd1854: data = 8'h7F;
            20'd1855: data = 8'h7F;
            20'd1856: data = 8'h7F;
            20'd1857: data = 8'h7F;
            20'd1858: data = 8'h80;
            20'd1859: data = 8'h80;
            20'd1860: data = 8'h7F;
            20'd1861: data = 8'h7F;
            20'd1862: data = 8'h80;
            20'd1863: data = 8'h80;
            20'd1864: data = 8'h7F;
            20'd1865: data = 8'h7F;
            20'd1866: data = 8'h80;
            20'd1867: data = 8'h80;
            20'd1868: data = 8'h7F;
            20'd1869: data = 8'h7F;
            20'd1870: data = 8'h80;
            20'd1871: data = 8'h80;
            20'd1872: data = 8'h7F;
            20'd1873: data = 8'h7F;
            20'd1874: data = 8'h7F;
            20'd1875: data = 8'h7F;
            20'd1876: data = 8'h7F;
            20'd1877: data = 8'h7F;
            20'd1878: data = 8'h80;
            20'd1879: data = 8'h80;
            20'd1880: data = 8'h7F;
            20'd1881: data = 8'h7F;
            20'd1882: data = 8'h7F;
            20'd1883: data = 8'h7F;
            20'd1884: data = 8'h7F;
            20'd1885: data = 8'h7F;
            20'd1886: data = 8'hA8;
            20'd1887: data = 8'hA8;
            20'd1888: data = 8'hAF;
            20'd1889: data = 8'hAF;
            20'd1890: data = 8'h9E;
            20'd1891: data = 8'h9E;
            20'd1892: data = 8'h8E;
            20'd1893: data = 8'h8E;
            20'd1894: data = 8'h82;
            20'd1895: data = 8'h82;
            20'd1896: data = 8'h77;
            20'd1897: data = 8'h77;
            20'd1898: data = 8'h6F;
            20'd1899: data = 8'h6F;
            20'd1900: data = 8'h6C;
            20'd1901: data = 8'h6C;
            20'd1902: data = 8'h6C;
            20'd1903: data = 8'h6C;
            20'd1904: data = 8'h21;
            20'd1905: data = 8'h21;
            20'd1906: data = 8'h3C;
            20'd1907: data = 8'h3C;
            20'd1908: data = 8'h51;
            20'd1909: data = 8'h51;
            20'd1910: data = 8'h65;
            20'd1911: data = 8'h65;
            20'd1912: data = 8'h76;
            20'd1913: data = 8'h76;
            20'd1914: data = 8'h84;
            20'd1915: data = 8'h84;
            20'd1916: data = 8'h8C;
            20'd1917: data = 8'h8C;
            20'd1918: data = 8'h94;
            20'd1919: data = 8'h94;
            20'd1920: data = 8'hE6;
            20'd1921: data = 8'hE6;
            20'd1922: data = 8'hCA;
            20'd1923: data = 8'hCA;
            20'd1924: data = 8'hB7;
            20'd1925: data = 8'hB7;
            20'd1926: data = 8'hA4;
            20'd1927: data = 8'hA4;
            20'd1928: data = 8'h94;
            20'd1929: data = 8'h94;
            20'd1930: data = 8'h86;
            20'd1931: data = 8'h86;
            20'd1932: data = 8'h7C;
            20'd1933: data = 8'h7C;
            20'd1934: data = 8'h74;
            20'd1935: data = 8'h74;
            20'd1936: data = 8'h1B;
            20'd1937: data = 8'h1B;
            20'd1938: data = 8'h38;
            20'd1939: data = 8'h38;
            20'd1940: data = 8'h4D;
            20'd1941: data = 8'h4D;
            20'd1942: data = 8'h60;
            20'd1943: data = 8'h60;
            20'd1944: data = 8'h70;
            20'd1945: data = 8'h70;
            20'd1946: data = 8'h7C;
            20'd1947: data = 8'h7C;
            20'd1948: data = 8'h86;
            20'd1949: data = 8'h86;
            20'd1950: data = 8'h91;
            20'd1951: data = 8'h91;
            20'd1952: data = 8'hE6;
            20'd1953: data = 8'hE6;
            20'd1954: data = 8'hCD;
            20'd1955: data = 8'hCD;
            20'd1956: data = 8'hB4;
            20'd1957: data = 8'hB4;
            20'd1958: data = 8'h9F;
            20'd1959: data = 8'h9F;
            20'd1960: data = 8'h8D;
            20'd1961: data = 8'h8D;
            20'd1962: data = 8'h80;
            20'd1963: data = 8'h80;
            20'd1964: data = 8'h74;
            20'd1965: data = 8'h74;
            20'd1966: data = 8'h6E;
            20'd1967: data = 8'h6E;
            20'd1968: data = 8'h24;
            20'd1969: data = 8'h24;
            20'd1970: data = 8'h2D;
            20'd1971: data = 8'h2D;
            20'd1972: data = 8'h42;
            20'd1973: data = 8'h42;
            20'd1974: data = 8'h58;
            20'd1975: data = 8'h58;
            20'd1976: data = 8'h6C;
            20'd1977: data = 8'h6C;
            20'd1978: data = 8'h7D;
            20'd1979: data = 8'h7D;
            20'd1980: data = 8'h89;
            20'd1981: data = 8'h89;
            20'd1982: data = 8'h92;
            20'd1983: data = 8'h92;
            20'd1984: data = 8'hBE;
            20'd1985: data = 8'hBE;
            20'd1986: data = 8'hD5;
            20'd1987: data = 8'hD5;
            20'd1988: data = 8'hC2;
            20'd1989: data = 8'hC2;
            20'd1990: data = 8'hAB;
            20'd1991: data = 8'hAB;
            20'd1992: data = 8'h99;
            20'd1993: data = 8'h99;
            20'd1994: data = 8'h87;
            20'd1995: data = 8'h87;
            20'd1996: data = 8'h7B;
            20'd1997: data = 8'h7B;
            20'd1998: data = 8'h70;
            20'd1999: data = 8'h70;
            20'd2000: data = 8'h60;
            20'd2001: data = 8'h60;
            20'd2002: data = 8'h28;
            20'd2003: data = 8'h28;
            20'd2004: data = 8'h3D;
            20'd2005: data = 8'h3D;
            20'd2006: data = 8'h53;
            20'd2007: data = 8'h53;
            20'd2008: data = 8'h65;
            20'd2009: data = 8'h65;
            20'd2010: data = 8'h77;
            20'd2011: data = 8'h77;
            20'd2012: data = 8'h83;
            20'd2013: data = 8'h83;
            20'd2014: data = 8'h8E;
            20'd2015: data = 8'h8E;
            20'd2016: data = 8'h8F;
            20'd2017: data = 8'h8F;
            20'd2018: data = 8'hDB;
            20'd2019: data = 8'hDB;
            20'd2020: data = 8'hC6;
            20'd2021: data = 8'hC6;
            20'd2022: data = 8'hAE;
            20'd2023: data = 8'hAE;
            20'd2024: data = 8'h9B;
            20'd2025: data = 8'h9B;
            20'd2026: data = 8'h88;
            20'd2027: data = 8'h88;
            20'd2028: data = 8'h7B;
            20'd2029: data = 8'h7B;
            20'd2030: data = 8'h72;
            20'd2031: data = 8'h72;
            20'd2032: data = 8'h6F;
            20'd2033: data = 8'h6F;
            20'd2034: data = 8'h1B;
            20'd2035: data = 8'h1B;
            20'd2036: data = 8'h36;
            20'd2037: data = 8'h36;
            20'd2038: data = 8'h4C;
            20'd2039: data = 8'h4C;
            20'd2040: data = 8'h62;
            20'd2041: data = 8'h62;
            20'd2042: data = 8'h74;
            20'd2043: data = 8'h74;
            20'd2044: data = 8'h82;
            20'd2045: data = 8'h82;
            20'd2046: data = 8'h8C;
            20'd2047: data = 8'h8C;
            20'd2048: data = 8'h95;
            20'd2049: data = 8'h95;
            20'd2050: data = 8'hEA;
            20'd2051: data = 8'hEA;
            20'd2052: data = 8'hCD;
            20'd2053: data = 8'hCD;
            20'd2054: data = 8'hB7;
            20'd2055: data = 8'hB7;
            20'd2056: data = 8'hA0;
            20'd2057: data = 8'hA0;
            20'd2058: data = 8'h8E;
            20'd2059: data = 8'h8E;
            20'd2060: data = 8'h7F;
            20'd2061: data = 8'h7F;
            20'd2062: data = 8'h75;
            20'd2063: data = 8'h75;
            20'd2064: data = 8'h6A;
            20'd2065: data = 8'h6A;
            20'd2066: data = 8'h14;
            20'd2067: data = 8'h14;
            20'd2068: data = 8'h31;
            20'd2069: data = 8'h31;
            20'd2070: data = 8'h47;
            20'd2071: data = 8'h47;
            20'd2072: data = 8'h5C;
            20'd2073: data = 8'h5C;
            20'd2074: data = 8'h6D;
            20'd2075: data = 8'h6D;
            20'd2076: data = 8'h7D;
            20'd2077: data = 8'h7D;
            20'd2078: data = 8'h89;
            20'd2079: data = 8'h89;
            20'd2080: data = 8'h90;
            20'd2081: data = 8'h90;
            20'd2082: data = 8'hDE;
            20'd2083: data = 8'hDE;
            20'd2084: data = 8'hD0;
            20'd2085: data = 8'hD0;
            20'd2086: data = 8'hBA;
            20'd2087: data = 8'hBA;
            20'd2088: data = 8'hA7;
            20'd2089: data = 8'hA7;
            20'd2090: data = 8'h93;
            20'd2091: data = 8'h93;
            20'd2092: data = 8'h82;
            20'd2093: data = 8'h82;
            20'd2094: data = 8'h77;
            20'd2095: data = 8'h77;
            20'd2096: data = 8'h70;
            20'd2097: data = 8'h70;
            20'd2098: data = 8'h3D;
            20'd2099: data = 8'h3D;
            20'd2100: data = 8'h2B;
            20'd2101: data = 8'h2B;
            20'd2102: data = 8'h40;
            20'd2103: data = 8'h40;
            20'd2104: data = 8'h54;
            20'd2105: data = 8'h54;
            20'd2106: data = 8'h69;
            20'd2107: data = 8'h69;
            20'd2108: data = 8'h79;
            20'd2109: data = 8'h79;
            20'd2110: data = 8'h86;
            20'd2111: data = 8'h86;
            20'd2112: data = 8'h90;
            20'd2113: data = 8'h90;
            20'd2114: data = 8'hA5;
            20'd2115: data = 8'hA5;
            20'd2116: data = 8'hD7;
            20'd2117: data = 8'hD7;
            20'd2118: data = 8'hC3;
            20'd2119: data = 8'hC3;
            20'd2120: data = 8'hAD;
            20'd2121: data = 8'hAD;
            20'd2122: data = 8'h99;
            20'd2123: data = 8'h99;
            20'd2124: data = 8'h89;
            20'd2125: data = 8'h89;
            20'd2126: data = 8'h7A;
            20'd2127: data = 8'h7A;
            20'd2128: data = 8'h70;
            20'd2129: data = 8'h70;
            20'd2130: data = 8'h6C;
            20'd2131: data = 8'h6C;
            20'd2132: data = 8'h23;
            20'd2133: data = 8'h23;
            20'd2134: data = 8'h3A;
            20'd2135: data = 8'h3A;
            20'd2136: data = 8'h50;
            20'd2137: data = 8'h50;
            20'd2138: data = 8'h63;
            20'd2139: data = 8'h63;
            20'd2140: data = 8'h74;
            20'd2141: data = 8'h74;
            20'd2142: data = 8'h83;
            20'd2143: data = 8'h83;
            20'd2144: data = 8'h8E;
            20'd2145: data = 8'h8E;
            20'd2146: data = 8'h92;
            20'd2147: data = 8'h92;
            20'd2148: data = 8'hE3;
            20'd2149: data = 8'hE3;
            20'd2150: data = 8'hC8;
            20'd2151: data = 8'hC8;
            20'd2152: data = 8'hB2;
            20'd2153: data = 8'hB2;
            20'd2154: data = 8'h9E;
            20'd2155: data = 8'h9E;
            20'd2156: data = 8'h8B;
            20'd2157: data = 8'h8B;
            20'd2158: data = 8'h7E;
            20'd2159: data = 8'h7E;
            20'd2160: data = 8'h74;
            20'd2161: data = 8'h74;
            20'd2162: data = 8'h6A;
            20'd2163: data = 8'h6A;
            20'd2164: data = 8'h15;
            20'd2165: data = 8'h15;
            20'd2166: data = 8'h33;
            20'd2167: data = 8'h33;
            20'd2168: data = 8'h4A;
            20'd2169: data = 8'h4A;
            20'd2170: data = 8'h60;
            20'd2171: data = 8'h60;
            20'd2172: data = 8'h71;
            20'd2173: data = 8'h71;
            20'd2174: data = 8'h7E;
            20'd2175: data = 8'h7E;
            20'd2176: data = 8'h8B;
            20'd2177: data = 8'h8B;
            20'd2178: data = 8'h94;
            20'd2179: data = 8'h94;
            20'd2180: data = 8'hEC;
            20'd2181: data = 8'hEC;
            20'd2182: data = 8'hCF;
            20'd2183: data = 8'hCF;
            20'd2184: data = 8'hB7;
            20'd2185: data = 8'hB7;
            20'd2186: data = 8'hA1;
            20'd2187: data = 8'hA1;
            20'd2188: data = 8'h92;
            20'd2189: data = 8'h92;
            20'd2190: data = 8'h81;
            20'd2191: data = 8'h81;
            20'd2192: data = 8'h75;
            20'd2193: data = 8'h75;
            20'd2194: data = 8'h6E;
            20'd2195: data = 8'h6E;
            20'd2196: data = 8'h1D;
            20'd2197: data = 8'h1D;
            20'd2198: data = 8'h2E;
            20'd2199: data = 8'h2E;
            20'd2200: data = 8'h45;
            20'd2201: data = 8'h45;
            20'd2202: data = 8'h5A;
            20'd2203: data = 8'h5A;
            20'd2204: data = 8'h6C;
            20'd2205: data = 8'h6C;
            20'd2206: data = 8'h7D;
            20'd2207: data = 8'h7D;
            20'd2208: data = 8'h87;
            20'd2209: data = 8'h87;
            20'd2210: data = 8'h90;
            20'd2211: data = 8'h90;
            20'd2212: data = 8'hC7;
            20'd2213: data = 8'hC7;
            20'd2214: data = 8'hD4;
            20'd2215: data = 8'hD4;
            20'd2216: data = 8'hBE;
            20'd2217: data = 8'hBE;
            20'd2218: data = 8'hA8;
            20'd2219: data = 8'hA8;
            20'd2220: data = 8'h93;
            20'd2221: data = 8'h93;
            20'd2222: data = 8'h86;
            20'd2223: data = 8'h86;
            20'd2224: data = 8'h7B;
            20'd2225: data = 8'h7B;
            20'd2226: data = 8'h70;
            20'd2227: data = 8'h70;
            20'd2228: data = 8'h57;
            20'd2229: data = 8'h57;
            20'd2230: data = 8'h28;
            20'd2231: data = 8'h28;
            20'd2232: data = 8'h3E;
            20'd2233: data = 8'h3E;
            20'd2234: data = 8'h54;
            20'd2235: data = 8'h54;
            20'd2236: data = 8'h68;
            20'd2237: data = 8'h68;
            20'd2238: data = 8'h77;
            20'd2239: data = 8'h77;
            20'd2240: data = 8'h84;
            20'd2241: data = 8'h84;
            20'd2242: data = 8'h8E;
            20'd2243: data = 8'h8E;
            20'd2244: data = 8'h94;
            20'd2245: data = 8'h94;
            20'd2246: data = 8'hDC;
            20'd2247: data = 8'hDC;
            20'd2248: data = 8'hC6;
            20'd2249: data = 8'hC6;
            20'd2250: data = 8'hB0;
            20'd2251: data = 8'hB0;
            20'd2252: data = 8'h9B;
            20'd2253: data = 8'h9B;
            20'd2254: data = 8'h89;
            20'd2255: data = 8'h89;
            20'd2256: data = 8'h7C;
            20'd2257: data = 8'h7C;
            20'd2258: data = 8'h72;
            20'd2259: data = 8'h72;
            20'd2260: data = 8'h6F;
            20'd2261: data = 8'h6F;
            20'd2262: data = 8'h1E;
            20'd2263: data = 8'h1E;
            20'd2264: data = 8'h36;
            20'd2265: data = 8'h36;
            20'd2266: data = 8'h4B;
            20'd2267: data = 8'h4B;
            20'd2268: data = 8'h61;
            20'd2269: data = 8'h61;
            20'd2270: data = 8'h74;
            20'd2271: data = 8'h74;
            20'd2272: data = 8'h82;
            20'd2273: data = 8'h82;
            20'd2274: data = 8'h8C;
            20'd2275: data = 8'h8C;
            20'd2276: data = 8'h93;
            20'd2277: data = 8'h93;
            20'd2278: data = 8'hE9;
            20'd2279: data = 8'hE9;
            20'd2280: data = 8'hCC;
            20'd2281: data = 8'hCC;
            20'd2282: data = 8'hB6;
            20'd2283: data = 8'hB6;
            20'd2284: data = 8'hA1;
            20'd2285: data = 8'hA1;
            20'd2286: data = 8'h8E;
            20'd2287: data = 8'h8E;
            20'd2288: data = 8'h7E;
            20'd2289: data = 8'h7E;
            20'd2290: data = 8'h74;
            20'd2291: data = 8'h74;
            20'd2292: data = 8'h6B;
            20'd2293: data = 8'h6B;
            20'd2294: data = 8'h13;
            20'd2295: data = 8'h13;
            20'd2296: data = 8'h30;
            20'd2297: data = 8'h30;
            20'd2298: data = 8'h48;
            20'd2299: data = 8'h48;
            20'd2300: data = 8'h5B;
            20'd2301: data = 8'h5B;
            20'd2302: data = 8'h6E;
            20'd2303: data = 8'h6E;
            20'd2304: data = 8'h7E;
            20'd2305: data = 8'h7E;
            20'd2306: data = 8'h8A;
            20'd2307: data = 8'h8A;
            20'd2308: data = 8'h92;
            20'd2309: data = 8'h92;
            20'd2310: data = 8'hE4;
            20'd2311: data = 8'hE4;
            20'd2312: data = 8'hD1;
            20'd2313: data = 8'hD1;
            20'd2314: data = 8'hBA;
            20'd2315: data = 8'hBA;
            20'd2316: data = 8'hA7;
            20'd2317: data = 8'hA7;
            20'd2318: data = 8'h94;
            20'd2319: data = 8'h94;
            20'd2320: data = 8'h84;
            20'd2321: data = 8'h84;
            20'd2322: data = 8'h77;
            20'd2323: data = 8'h77;
            20'd2324: data = 8'h6F;
            20'd2325: data = 8'h6F;
            20'd2326: data = 8'h32;
            20'd2327: data = 8'h32;
            20'd2328: data = 8'h2C;
            20'd2329: data = 8'h2C;
            20'd2330: data = 8'h41;
            20'd2331: data = 8'h41;
            20'd2332: data = 8'h55;
            20'd2333: data = 8'h55;
            20'd2334: data = 8'h69;
            20'd2335: data = 8'h69;
            20'd2336: data = 8'h79;
            20'd2337: data = 8'h79;
            20'd2338: data = 8'h87;
            20'd2339: data = 8'h87;
            20'd2340: data = 8'h91;
            20'd2341: data = 8'h91;
            20'd2342: data = 8'hAE;
            20'd2343: data = 8'hAE;
            20'd2344: data = 8'hD6;
            20'd2345: data = 8'hD6;
            20'd2346: data = 8'hC1;
            20'd2347: data = 8'hC1;
            20'd2348: data = 8'hAB;
            20'd2349: data = 8'hAB;
            20'd2350: data = 8'h98;
            20'd2351: data = 8'h98;
            20'd2352: data = 8'h89;
            20'd2353: data = 8'h89;
            20'd2354: data = 8'h7A;
            20'd2355: data = 8'h7A;
            20'd2356: data = 8'h6F;
            20'd2357: data = 8'h6F;
            20'd2358: data = 8'h67;
            20'd2359: data = 8'h67;
            20'd2360: data = 8'h24;
            20'd2361: data = 8'h24;
            20'd2362: data = 8'h3B;
            20'd2363: data = 8'h3B;
            20'd2364: data = 8'h53;
            20'd2365: data = 8'h53;
            20'd2366: data = 8'h66;
            20'd2367: data = 8'h66;
            20'd2368: data = 8'h74;
            20'd2369: data = 8'h74;
            20'd2370: data = 8'h82;
            20'd2371: data = 8'h82;
            20'd2372: data = 8'h8C;
            20'd2373: data = 8'h8C;
            20'd2374: data = 8'h8F;
            20'd2375: data = 8'h90;
            20'd2376: data = 8'hE0;
            20'd2377: data = 8'hE0;
            20'd2378: data = 8'hC8;
            20'd2379: data = 8'hC8;
            20'd2380: data = 8'hB0;
            20'd2381: data = 8'hB0;
            20'd2382: data = 8'h9D;
            20'd2383: data = 8'h9D;
            20'd2384: data = 8'h8C;
            20'd2385: data = 8'h8C;
            20'd2386: data = 8'h7F;
            20'd2387: data = 8'h7F;
            20'd2388: data = 8'h74;
            20'd2389: data = 8'h74;
            20'd2390: data = 8'h6C;
            20'd2391: data = 8'h6C;
            20'd2392: data = 8'h18;
            20'd2393: data = 8'h18;
            20'd2394: data = 8'h34;
            20'd2395: data = 8'h34;
            20'd2396: data = 8'h4A;
            20'd2397: data = 8'h4A;
            20'd2398: data = 8'h5F;
            20'd2399: data = 8'h5F;
            20'd2400: data = 8'h72;
            20'd2401: data = 8'h72;
            20'd2402: data = 8'h7F;
            20'd2403: data = 8'h7F;
            20'd2404: data = 8'h8A;
            20'd2405: data = 8'h8A;
            20'd2406: data = 8'h96;
            20'd2407: data = 8'h96;
            20'd2408: data = 8'hED;
            20'd2409: data = 8'hED;
            20'd2410: data = 8'hCF;
            20'd2411: data = 8'hCF;
            20'd2412: data = 8'hB7;
            20'd2413: data = 8'hB7;
            20'd2414: data = 8'hA3;
            20'd2415: data = 8'hA3;
            20'd2416: data = 8'h8F;
            20'd2417: data = 8'h8F;
            20'd2418: data = 8'h81;
            20'd2419: data = 8'h81;
            20'd2420: data = 8'h74;
            20'd2421: data = 8'h74;
            20'd2422: data = 8'h6C;
            20'd2423: data = 8'h6C;
            20'd2424: data = 8'h16;
            20'd2425: data = 8'h16;
            20'd2426: data = 8'h2F;
            20'd2427: data = 8'h2F;
            20'd2428: data = 8'h46;
            20'd2429: data = 8'h46;
            20'd2430: data = 8'h5A;
            20'd2431: data = 8'h5A;
            20'd2432: data = 8'h6D;
            20'd2433: data = 8'h6D;
            20'd2434: data = 8'h7D;
            20'd2435: data = 8'h7D;
            20'd2436: data = 8'h89;
            20'd2437: data = 8'h89;
            20'd2438: data = 8'h90;
            20'd2439: data = 8'h90;
            20'd2440: data = 8'hD3;
            20'd2441: data = 8'hD3;
            20'd2442: data = 8'hD1;
            20'd2443: data = 8'hD1;
            20'd2444: data = 8'hBD;
            20'd2445: data = 8'hBD;
            20'd2446: data = 8'hA7;
            20'd2447: data = 8'hA7;
            20'd2448: data = 8'h95;
            20'd2449: data = 8'h95;
            20'd2450: data = 8'h84;
            20'd2451: data = 8'h84;
            20'd2452: data = 8'h78;
            20'd2453: data = 8'h78;
            20'd2454: data = 8'h70;
            20'd2455: data = 8'h70;
            20'd2456: data = 8'h4C;
            20'd2457: data = 8'h4C;
            20'd2458: data = 8'h2A;
            20'd2459: data = 8'h2A;
            20'd2460: data = 8'h3F;
            20'd2461: data = 8'h3F;
            20'd2462: data = 8'h55;
            20'd2463: data = 8'h55;
            20'd2464: data = 8'h69;
            20'd2465: data = 8'h69;
            20'd2466: data = 8'h78;
            20'd2467: data = 8'h78;
            20'd2468: data = 8'h86;
            20'd2469: data = 8'h86;
            20'd2470: data = 8'h8F;
            20'd2471: data = 8'h8F;
            20'd2472: data = 8'h9B;
            20'd2473: data = 8'h9B;
            20'd2474: data = 8'hDB;
            20'd2475: data = 8'hDB;
            20'd2476: data = 8'hC3;
            20'd2477: data = 8'hC3;
            20'd2478: data = 8'hAC;
            20'd2479: data = 8'hAC;
            20'd2480: data = 8'h9A;
            20'd2481: data = 8'h9A;
            20'd2482: data = 8'h89;
            20'd2483: data = 8'h89;
            20'd2484: data = 8'h7A;
            20'd2485: data = 8'h7A;
            20'd2486: data = 8'h71;
            20'd2487: data = 8'h71;
            20'd2488: data = 8'h6E;
            20'd2489: data = 8'h6E;
            20'd2490: data = 8'h21;
            20'd2491: data = 8'h21;
            20'd2492: data = 8'h3A;
            20'd2493: data = 8'h3A;
            20'd2494: data = 8'h4F;
            20'd2495: data = 8'h4F;
            20'd2496: data = 8'h62;
            20'd2497: data = 8'h62;
            20'd2498: data = 8'h75;
            20'd2499: data = 8'h75;
            20'd2500: data = 8'h83;
            20'd2501: data = 8'h83;
            20'd2502: data = 8'h8C;
            20'd2503: data = 8'h8C;
            20'd2504: data = 8'h92;
            20'd2505: data = 8'h92;
            20'd2506: data = 8'hE6;
            20'd2507: data = 8'hE6;
            20'd2508: data = 8'hC9;
            20'd2509: data = 8'hC9;
            20'd2510: data = 8'hB4;
            20'd2511: data = 8'hB4;
            20'd2512: data = 8'hA0;
            20'd2513: data = 8'hA0;
            20'd2514: data = 8'h8D;
            20'd2515: data = 8'h8D;
            20'd2516: data = 8'h7F;
            20'd2517: data = 8'h7F;
            20'd2518: data = 8'h75;
            20'd2519: data = 8'h75;
            20'd2520: data = 8'h6A;
            20'd2521: data = 8'h6A;
            20'd2522: data = 8'h13;
            20'd2523: data = 8'h13;
            20'd2524: data = 8'h31;
            20'd2525: data = 8'h31;
            20'd2526: data = 8'h58;
            20'd2527: data = 8'h58;
            20'd2528: data = 8'h67;
            20'd2529: data = 8'h67;
            20'd2530: data = 8'h75;
            20'd2531: data = 8'h75;
            20'd2532: data = 8'h80;
            20'd2533: data = 8'h80;
            20'd2534: data = 8'h8A;
            20'd2535: data = 8'h8A;
            20'd2536: data = 8'h91;
            20'd2537: data = 8'h91;
            20'd2538: data = 8'h93;
            20'd2539: data = 8'h93;
            20'd2540: data = 8'h94;
            20'd2541: data = 8'h94;
            20'd2542: data = 8'h93;
            20'd2543: data = 8'h93;
            20'd2544: data = 8'h92;
            20'd2545: data = 8'h92;
            20'd2546: data = 8'h8C;
            20'd2547: data = 8'h8C;
            20'd2548: data = 8'h89;
            20'd2549: data = 8'h89;
            20'd2550: data = 8'h85;
            20'd2551: data = 8'h85;
            20'd2552: data = 8'h82;
            20'd2553: data = 8'h82;
            20'd2554: data = 8'h82;
            20'd2555: data = 8'h82;
            20'd2556: data = 8'h80;
            20'd2557: data = 8'h80;
            20'd2558: data = 8'h81;
            20'd2559: data = 8'h81;
            20'd2560: data = 8'h82;
            20'd2561: data = 8'h82;
            20'd2562: data = 8'h83;
            20'd2563: data = 8'h83;
            20'd2564: data = 8'h83;
            20'd2565: data = 8'h83;
            20'd2566: data = 8'h83;
            20'd2567: data = 8'h83;
            20'd2568: data = 8'h82;
            20'd2569: data = 8'h82;
            20'd2570: data = 8'h83;
            20'd2571: data = 8'h83;
            20'd2572: data = 8'h82;
            20'd2573: data = 8'h82;
            20'd2574: data = 8'h80;
            20'd2575: data = 8'h80;
            20'd2576: data = 8'h7D;
            20'd2577: data = 8'h7D;
            20'd2578: data = 8'h7B;
            20'd2579: data = 8'h7B;
            20'd2580: data = 8'h7A;
            20'd2581: data = 8'h7A;
            20'd2582: data = 8'h79;
            20'd2583: data = 8'h79;
            20'd2584: data = 8'h78;
            20'd2585: data = 8'h78;
            20'd2586: data = 8'h78;
            20'd2587: data = 8'h78;
            20'd2588: data = 8'h79;
            20'd2589: data = 8'h79;
            20'd2590: data = 8'h79;
            20'd2591: data = 8'h79;
            20'd2592: data = 8'h7B;
            20'd2593: data = 8'h7B;
            20'd2594: data = 8'h7B;
            20'd2595: data = 8'h7B;
            20'd2596: data = 8'h7D;
            20'd2597: data = 8'h7D;
            20'd2598: data = 8'h80;
            20'd2599: data = 8'h80;
            20'd2600: data = 8'h81;
            20'd2601: data = 8'h81;
            20'd2602: data = 8'h82;
            20'd2603: data = 8'h82;
            20'd2604: data = 8'h82;
            20'd2605: data = 8'h82;
            20'd2606: data = 8'h84;
            20'd2607: data = 8'h84;
            20'd2608: data = 8'h83;
            20'd2609: data = 8'h83;
            20'd2610: data = 8'h82;
            20'd2611: data = 8'h82;
            20'd2612: data = 8'h83;
            20'd2613: data = 8'h83;
            20'd2614: data = 8'h82;
            20'd2615: data = 8'h82;
            20'd2616: data = 8'h80;
            20'd2617: data = 8'h80;
            20'd2618: data = 8'h80;
            20'd2619: data = 8'h80;
            20'd2620: data = 8'h80;
            20'd2621: data = 8'h80;
            20'd2622: data = 8'h7F;
            20'd2623: data = 8'h7F;
            20'd2624: data = 8'h7E;
            20'd2625: data = 8'h7E;
            20'd2626: data = 8'h80;
            20'd2627: data = 8'h80;
            20'd2628: data = 8'h7F;
            20'd2629: data = 8'h7F;
            20'd2630: data = 8'h7F;
            20'd2631: data = 8'h7F;
            20'd2632: data = 8'h80;
            20'd2633: data = 8'h80;
            20'd2634: data = 8'h7F;
            20'd2635: data = 8'h7F;
            20'd2636: data = 8'h7F;
            20'd2637: data = 8'h7F;
            20'd2638: data = 8'h7F;
            20'd2639: data = 8'h7F;
            20'd2640: data = 8'h7F;
            20'd2641: data = 8'h7F;
            20'd2642: data = 8'h7E;
            20'd2643: data = 8'h7E;
            20'd2644: data = 8'h7E;
            20'd2645: data = 8'h7E;
            20'd2646: data = 8'h7F;
            20'd2647: data = 8'h7F;
            20'd2648: data = 8'h7E;
            20'd2649: data = 8'h7E;
            20'd2650: data = 8'h7E;
            20'd2651: data = 8'h7E;
            20'd2652: data = 8'h7E;
            20'd2653: data = 8'h7E;
            20'd2654: data = 8'h7F;
            20'd2655: data = 8'h7F;
            20'd2656: data = 8'h7F;
            20'd2657: data = 8'h7F;
            20'd2658: data = 8'h7F;
            20'd2659: data = 8'h7F;
            20'd2660: data = 8'h7F;
            20'd2661: data = 8'h7F;
            20'd2662: data = 8'h80;
            20'd2663: data = 8'h80;
            20'd2664: data = 8'h80;
            20'd2665: data = 8'h80;
            20'd2666: data = 8'h80;
            20'd2667: data = 8'h80;
            20'd2668: data = 8'h80;
            20'd2669: data = 8'h80;
            20'd2670: data = 8'h80;
            20'd2671: data = 8'h80;
            20'd2672: data = 8'h80;
            20'd2673: data = 8'h80;
            20'd2674: data = 8'h80;
            20'd2675: data = 8'h80;
            20'd2676: data = 8'h80;
            20'd2677: data = 8'h80;
            20'd2678: data = 8'h80;
            20'd2679: data = 8'h80;
            20'd2680: data = 8'h80;
            20'd2681: data = 8'h80;
            20'd2682: data = 8'h80;
            20'd2683: data = 8'h80;
            20'd2684: data = 8'h80;
            20'd2685: data = 8'h80;
            20'd2686: data = 8'h80;
            20'd2687: data = 8'h80;
            20'd2688: data = 8'h80;
            20'd2689: data = 8'h80;
            20'd2690: data = 8'h80;
            20'd2691: data = 8'h80;
            20'd2692: data = 8'h80;
            20'd2693: data = 8'h80;
            20'd2694: data = 8'h7F;
            20'd2695: data = 8'h7F;
            20'd2696: data = 8'h7F;
            20'd2697: data = 8'h7F;
            20'd2698: data = 8'h7F;
            20'd2699: data = 8'h7F;
            20'd2700: data = 8'h7F;
            20'd2701: data = 8'h7F;
            20'd2702: data = 8'h7F;
            20'd2703: data = 8'h7F;
            20'd2704: data = 8'h7F;
            20'd2705: data = 8'h7F;
            20'd2706: data = 8'h7F;
            20'd2707: data = 8'h7F;
            20'd2708: data = 8'h7F;
            20'd2709: data = 8'h7F;
            20'd2710: data = 8'h7F;
            20'd2711: data = 8'h7F;
            20'd2712: data = 8'h7F;
            20'd2713: data = 8'h7F;
            20'd2714: data = 8'h7F;
            20'd2715: data = 8'h7F;
            20'd2716: data = 8'h7F;
            20'd2717: data = 8'h7F;
            20'd2718: data = 8'h7F;
            20'd2719: data = 8'h7F;
            20'd2720: data = 8'h7F;
            20'd2721: data = 8'h7F;
            20'd2722: data = 8'h7F;
            20'd2723: data = 8'h7F;
            20'd2724: data = 8'h7F;
            20'd2725: data = 8'h7F;
            20'd2726: data = 8'h7F;
            20'd2727: data = 8'h7F;
            20'd2728: data = 8'h7F;
            20'd2729: data = 8'h7F;
            20'd2730: data = 8'h7F;
            20'd2731: data = 8'h80;
            20'd2732: data = 8'h80;
            20'd2733: data = 8'h80;
            20'd2734: data = 8'h80;
            20'd2735: data = 8'h80;
            20'd2736: data = 8'h80;
            20'd2737: data = 8'h80;
            20'd2738: data = 8'h80;
            20'd2739: data = 8'h80;
            20'd2740: data = 8'h80;
            20'd2741: data = 8'h80;
            20'd2742: data = 8'h80;
            20'd2743: data = 8'h80;
            20'd2744: data = 8'h80;
            20'd2745: data = 8'h80;
            20'd2746: data = 8'h80;
            20'd2747: data = 8'h80;
            20'd2748: data = 8'h80;
            20'd2749: data = 8'h80;
            20'd2750: data = 8'h80;
            20'd2751: data = 8'h80;
            20'd2752: data = 8'h80;
            20'd2753: data = 8'h80;
            20'd2754: data = 8'h80;
            20'd2755: data = 8'h80;
            20'd2756: data = 8'h80;
            20'd2757: data = 8'h80;
            20'd2758: data = 8'h80;
            20'd2759: data = 8'h7F;
            20'd2760: data = 8'h80;
            20'd2761: data = 8'h7F;
            20'd2762: data = 8'h7F;
            20'd2763: data = 8'h7F;
            20'd2764: data = 8'h7F;
            20'd2765: data = 8'h7F;
            20'd2766: data = 8'h7F;
            20'd2767: data = 8'h7F;
            20'd2768: data = 8'h7F;
            20'd2769: data = 8'h7F;
            20'd2770: data = 8'h7F;
            20'd2771: data = 8'h7F;
            20'd2772: data = 8'h7F;
            20'd2773: data = 8'h7F;
            20'd2774: data = 8'h7F;
            20'd2775: data = 8'h7F;
            20'd2776: data = 8'h80;
            20'd2777: data = 8'h7F;
            20'd2778: data = 8'h7F;
            20'd2779: data = 8'h7F;
            20'd2780: data = 8'h7F;
            20'd2781: data = 8'h7F;
            20'd2782: data = 8'h7F;
            20'd2783: data = 8'h7F;
            20'd2784: data = 8'h7F;
            20'd2785: data = 8'h7F;
            20'd2786: data = 8'h7F;
            20'd2787: data = 8'h7F;
            20'd2788: data = 8'h7F;
            20'd2789: data = 8'h80;
            20'd2790: data = 8'h80;
            20'd2791: data = 8'h80;
            20'd2792: data = 8'h7F;
            20'd2793: data = 8'h7F;
            20'd2794: data = 8'h80;
            20'd2795: data = 8'h7F;
            20'd2796: data = 8'h80;
            20'd2797: data = 8'h80;
            20'd2798: data = 8'h80;
            20'd2799: data = 8'h80;
            20'd2800: data = 8'h80;
            20'd2801: data = 8'h80;
            20'd2802: data = 8'h80;
            20'd2803: data = 8'h80;
            20'd2804: data = 8'h80;
            20'd2805: data = 8'h80;
            20'd2806: data = 8'h80;
            20'd2807: data = 8'h80;
            20'd2808: data = 8'h80;
            20'd2809: data = 8'h80;
            20'd2810: data = 8'h80;
            20'd2811: data = 8'h80;
            20'd2812: data = 8'h80;
            20'd2813: data = 8'h80;
            20'd2814: data = 8'h80;
            20'd2815: data = 8'h80;
            20'd2816: data = 8'h7F;
            20'd2817: data = 8'h7F;
            20'd2818: data = 8'h7F;
            20'd2819: data = 8'h7F;
            20'd2820: data = 8'h80;
            20'd2821: data = 8'h80;
            20'd2822: data = 8'h80;
            20'd2823: data = 8'h80;
            20'd2824: data = 8'h80;
            20'd2825: data = 8'h7F;
            20'd2826: data = 8'h80;
            20'd2827: data = 8'h7F;
            20'd2828: data = 8'h80;
            20'd2829: data = 8'h7F;
            20'd2830: data = 8'h7F;
            20'd2831: data = 8'h80;
            20'd2832: data = 8'h80;
            20'd2833: data = 8'h80;
            20'd2834: data = 8'h7F;
            20'd2835: data = 8'h7F;
            20'd2836: data = 8'h7F;
            20'd2837: data = 8'h7F;
            20'd2838: data = 8'h80;
            20'd2839: data = 8'h7F;
            20'd2840: data = 8'h7F;
            20'd2841: data = 8'h80;
            20'd2842: data = 8'h80;
            20'd2843: data = 8'h7F;
            20'd2844: data = 8'h7F;
            20'd2845: data = 8'h80;
            20'd2846: data = 8'h80;
            20'd2847: data = 8'h7F;
            20'd2848: data = 8'h7F;
            20'd2849: data = 8'h80;
            20'd2850: data = 8'h7F;
            20'd2851: data = 8'h7F;
            20'd2852: data = 8'h7F;
            20'd2853: data = 8'h80;
            20'd2854: data = 8'h7F;
            20'd2855: data = 8'h7F;
            20'd2856: data = 8'h7F;
            20'd2857: data = 8'h7F;
            20'd2858: data = 8'h80;
            20'd2859: data = 8'h7F;
            20'd2860: data = 8'h7F;
            20'd2861: data = 8'h7F;
            20'd2862: data = 8'h7F;
            20'd2863: data = 8'h7F;
            20'd2864: data = 8'h7F;
            20'd2865: data = 8'h80;
            20'd2866: data = 8'h7F;
            20'd2867: data = 8'h7F;
            20'd2868: data = 8'h7F;
            20'd2869: data = 8'h7F;
            20'd2870: data = 8'h7F;
            20'd2871: data = 8'h80;
            20'd2872: data = 8'h80;
            20'd2873: data = 8'h80;
            20'd2874: data = 8'h80;
            20'd2875: data = 8'h80;
            20'd2876: data = 8'h7F;
            20'd2877: data = 8'h7F;
            20'd2878: data = 8'h7F;
            20'd2879: data = 8'h80;
            20'd2880: data = 8'h80;
            20'd2881: data = 8'h7F;
            20'd2882: data = 8'h80;
            20'd2883: data = 8'h7F;
            20'd2884: data = 8'h7F;
            20'd2885: data = 8'h7F;
            20'd2886: data = 8'h7F;
            20'd2887: data = 8'h80;
            20'd2888: data = 8'h80;
            20'd2889: data = 8'h7F;
            20'd2890: data = 8'h7F;
            20'd2891: data = 8'h80;
            20'd2892: data = 8'h80;
            20'd2893: data = 8'h80;
            20'd2894: data = 8'h7F;
            20'd2895: data = 8'h80;
            20'd2896: data = 8'h80;
            20'd2897: data = 8'h7F;
            20'd2898: data = 8'h80;
            20'd2899: data = 8'h80;
            20'd2900: data = 8'h80;
            20'd2901: data = 8'h7F;
            20'd2902: data = 8'h80;
            20'd2903: data = 8'h80;
            20'd2904: data = 8'h80;
            20'd2905: data = 8'h7F;
            20'd2906: data = 8'h7F;
            20'd2907: data = 8'h7F;
            20'd2908: data = 8'h80;
            20'd2909: data = 8'h80;
            20'd2910: data = 8'h80;
            20'd2911: data = 8'h80;
            20'd2912: data = 8'h80;
            20'd2913: data = 8'h80;
            20'd2914: data = 8'h7F;
            20'd2915: data = 8'h7F;
            20'd2916: data = 8'h80;
            20'd2917: data = 8'h80;
            20'd2918: data = 8'h80;
            20'd2919: data = 8'h80;
            20'd2920: data = 8'h7F;
            20'd2921: data = 8'h80;
            20'd2922: data = 8'h7F;
            20'd2923: data = 8'h80;
            20'd2924: data = 8'h80;
            20'd2925: data = 8'h80;
            20'd2926: data = 8'h7F;
            20'd2927: data = 8'h80;
            20'd2928: data = 8'h80;
            20'd2929: data = 8'h7F;
            20'd2930: data = 8'h7F;
            20'd2931: data = 8'h7F;
            20'd2932: data = 8'h7F;
            20'd2933: data = 8'h7F;
            20'd2934: data = 8'h7F;
            20'd2935: data = 8'h80;
            20'd2936: data = 8'h80;
            20'd2937: data = 8'h80;
            20'd2938: data = 8'h7F;
            20'd2939: data = 8'h7F;
            20'd2940: data = 8'h7F;
            20'd2941: data = 8'h7F;
            20'd2942: data = 8'h7F;
            20'd2943: data = 8'h7F;
            20'd2944: data = 8'h7F;
            20'd2945: data = 8'h7F;
            20'd2946: data = 8'h7F;
            20'd2947: data = 8'h80;
            20'd2948: data = 8'h80;
            20'd2949: data = 8'h7F;
            20'd2950: data = 8'h7F;
            20'd2951: data = 8'h7F;
            20'd2952: data = 8'h80;
            20'd2953: data = 8'h7F;
            20'd2954: data = 8'h80;
            20'd2955: data = 8'h80;
            20'd2956: data = 8'h7F;
            20'd2957: data = 8'h7F;
            20'd2958: data = 8'h7F;
            20'd2959: data = 8'h7F;
            20'd2960: data = 8'h7F;
            20'd2961: data = 8'h7F;
            20'd2962: data = 8'h80;
            20'd2963: data = 8'h7F;
            20'd2964: data = 8'h7F;
            20'd2965: data = 8'h7F;
            20'd2966: data = 8'h80;
            20'd2967: data = 8'h80;
            20'd2968: data = 8'h80;
            20'd2969: data = 8'h80;
            20'd2970: data = 8'h80;
            20'd2971: data = 8'h7F;
            20'd2972: data = 8'h7F;
            20'd2973: data = 8'h7F;
            20'd2974: data = 8'h80;
            20'd2975: data = 8'h80;
            20'd2976: data = 8'h80;
            20'd2977: data = 8'h80;
            20'd2978: data = 8'h7F;
            20'd2979: data = 8'h80;
            20'd2980: data = 8'h80;
            20'd2981: data = 8'h80;
            20'd2982: data = 8'h80;
            20'd2983: data = 8'h7F;
            20'd2984: data = 8'h80;
            20'd2985: data = 8'h80;
            20'd2986: data = 8'h7F;
            20'd2987: data = 8'h7F;
            20'd2988: data = 8'h7F;
            20'd2989: data = 8'h80;
            20'd2990: data = 8'h80;
            20'd2991: data = 8'h7F;
            20'd2992: data = 8'h80;
            20'd2993: data = 8'h80;
            20'd2994: data = 8'h80;
            20'd2995: data = 8'h80;
            20'd2996: data = 8'h80;
            20'd2997: data = 8'h80;
            20'd2998: data = 8'h7F;
            20'd2999: data = 8'h7F;
            20'd3000: data = 8'h80;
            20'd3001: data = 8'h80;
            20'd3002: data = 8'h80;
            20'd3003: data = 8'h7F;
            20'd3004: data = 8'h7F;
            20'd3005: data = 8'h80;
            20'd3006: data = 8'h80;
            20'd3007: data = 8'h80;
            20'd3008: data = 8'h80;
            20'd3009: data = 8'h80;
            20'd3010: data = 8'h7F;
            20'd3011: data = 8'h80;
            20'd3012: data = 8'h7F;
            20'd3013: data = 8'h7F;
            20'd3014: data = 8'h80;
            20'd3015: data = 8'h80;
            20'd3016: data = 8'h7F;
            20'd3017: data = 8'h80;
            20'd3018: data = 8'h80;
            20'd3019: data = 8'h80;
            20'd3020: data = 8'h80;
            20'd3021: data = 8'h7F;
            20'd3022: data = 8'h80;
            20'd3023: data = 8'h80;
            20'd3024: data = 8'h80;
            20'd3025: data = 8'h80;
            20'd3026: data = 8'h80;
            20'd3027: data = 8'h80;
            20'd3028: data = 8'h80;
            20'd3029: data = 8'h80;
            20'd3030: data = 8'h80;
            20'd3031: data = 8'h80;
            20'd3032: data = 8'h7F;
            20'd3033: data = 8'h80;
            20'd3034: data = 8'h80;
            20'd3035: data = 8'h7F;
            20'd3036: data = 8'h80;
            20'd3037: data = 8'h7F;
            20'd3038: data = 8'h7F;
            20'd3039: data = 8'h7F;
            20'd3040: data = 8'h80;
            20'd3041: data = 8'h80;
            20'd3042: data = 8'h80;
            20'd3043: data = 8'h80;
            20'd3044: data = 8'h7F;
            20'd3045: data = 8'h80;
            20'd3046: data = 8'h80;
            20'd3047: data = 8'h80;
            20'd3048: data = 8'h80;
            20'd3049: data = 8'h80;
            20'd3050: data = 8'h7F;
            20'd3051: data = 8'h80;
            20'd3052: data = 8'h7F;
            20'd3053: data = 8'h7F;
            20'd3054: data = 8'h7F;
            20'd3055: data = 8'h7F;
            20'd3056: data = 8'h7F;
            20'd3057: data = 8'h7F;
            20'd3058: data = 8'h80;
            20'd3059: data = 8'h7F;
            20'd3060: data = 8'h80;
            20'd3061: data = 8'h7F;
            20'd3062: data = 8'h7F;
            20'd3063: data = 8'h80;
            20'd3064: data = 8'h80;
            20'd3065: data = 8'h80;
            20'd3066: data = 8'h7F;
            20'd3067: data = 8'h7F;
            20'd3068: data = 8'h7F;
            20'd3069: data = 8'h80;
            20'd3070: data = 8'h7F;
            20'd3071: data = 8'h80;
            20'd3072: data = 8'h80;
            20'd3073: data = 8'h80;
            20'd3074: data = 8'h7F;
            20'd3075: data = 8'h7F;
            20'd3076: data = 8'h7F;
            20'd3077: data = 8'h7F;
            20'd3078: data = 8'h7F;
            20'd3079: data = 8'h80;
            20'd3080: data = 8'h80;
            20'd3081: data = 8'h80;
            20'd3082: data = 8'h7F;
            20'd3083: data = 8'h7F;
            20'd3084: data = 8'h80;
            20'd3085: data = 8'h7F;
            20'd3086: data = 8'h7F;
            20'd3087: data = 8'h80;
            20'd3088: data = 8'h7F;
            20'd3089: data = 8'h7F;
            20'd3090: data = 8'h7F;
            20'd3091: data = 8'h7F;
            20'd3092: data = 8'h7F;
            20'd3093: data = 8'h7F;
            20'd3094: data = 8'h7F;
            20'd3095: data = 8'h7F;
            20'd3096: data = 8'h7F;
            20'd3097: data = 8'h7F;
            20'd3098: data = 8'h7F;
            20'd3099: data = 8'h7F;
            20'd3100: data = 8'h80;
            20'd3101: data = 8'h80;
            20'd3102: data = 8'h7F;
            20'd3103: data = 8'h7F;
            20'd3104: data = 8'h80;
            20'd3105: data = 8'h80;
            20'd3106: data = 8'h7F;
            20'd3107: data = 8'h80;
            20'd3108: data = 8'h80;
            20'd3109: data = 8'h7F;
            20'd3110: data = 8'h80;
            20'd3111: data = 8'h80;
            20'd3112: data = 8'h80;
            20'd3113: data = 8'h80;
            20'd3114: data = 8'h7F;
            20'd3115: data = 8'h80;
            20'd3116: data = 8'h80;
            20'd3117: data = 8'h80;
            20'd3118: data = 8'h80;
            20'd3119: data = 8'h80;
            20'd3120: data = 8'h80;
            20'd3121: data = 8'h7F;
            20'd3122: data = 8'h80;
            20'd3123: data = 8'h80;
            20'd3124: data = 8'h80;
            20'd3125: data = 8'h7F;
            20'd3126: data = 8'h7F;
            20'd3127: data = 8'h7F;
            20'd3128: data = 8'h80;
            20'd3129: data = 8'h80;
            20'd3130: data = 8'h80;
            20'd3131: data = 8'h7F;
            20'd3132: data = 8'h80;
            20'd3133: data = 8'h80;
            20'd3134: data = 8'h7F;
            20'd3135: data = 8'h7F;
            20'd3136: data = 8'h80;
            20'd3137: data = 8'h7F;
            20'd3138: data = 8'h80;
            20'd3139: data = 8'h80;
            20'd3140: data = 8'h7F;
            20'd3141: data = 8'h7F;
            20'd3142: data = 8'h80;
            20'd3143: data = 8'h7F;
            20'd3144: data = 8'h7F;
            20'd3145: data = 8'h7F;
            20'd3146: data = 8'h7F;
            20'd3147: data = 8'h7F;
            20'd3148: data = 8'h80;
            20'd3149: data = 8'h7F;
            20'd3150: data = 8'h7F;
            20'd3151: data = 8'h7F;
            20'd3152: data = 8'h80;
            20'd3153: data = 8'h80;
            20'd3154: data = 8'h7F;
            20'd3155: data = 8'h7F;
            20'd3156: data = 8'h7F;
            20'd3157: data = 8'h80;
            20'd3158: data = 8'h80;
            20'd3159: data = 8'h80;
            20'd3160: data = 8'h7F;
            20'd3161: data = 8'h7F;
            20'd3162: data = 8'h7F;
            20'd3163: data = 8'h7F;
            20'd3164: data = 8'h80;
            20'd3165: data = 8'h7F;
            20'd3166: data = 8'h7F;
            20'd3167: data = 8'h80;
            20'd3168: data = 8'h80;
            20'd3169: data = 8'h7F;
            20'd3170: data = 8'h80;
            20'd3171: data = 8'h80;
            20'd3172: data = 8'h80;
            20'd3173: data = 8'h7F;
            20'd3174: data = 8'h80;
            20'd3175: data = 8'h80;
            20'd3176: data = 8'h80;
            20'd3177: data = 8'h80;
            20'd3178: data = 8'h80;
            20'd3179: data = 8'h7F;
            20'd3180: data = 8'h7F;
            20'd3181: data = 8'h80;
            20'd3182: data = 8'h80;
            20'd3183: data = 8'h80;
            20'd3184: data = 8'h7F;
            20'd3185: data = 8'h80;
            20'd3186: data = 8'h80;
            20'd3187: data = 8'h7F;
            20'd3188: data = 8'h7F;
            20'd3189: data = 8'h80;
            20'd3190: data = 8'h7F;
            20'd3191: data = 8'h80;
            20'd3192: data = 8'h80;
            20'd3193: data = 8'h7F;
            20'd3194: data = 8'h7F;
            20'd3195: data = 8'h7F;
            20'd3196: data = 8'h80;
            20'd3197: data = 8'h7F;
            20'd3198: data = 8'h80;
            20'd3199: data = 8'h80;
            20'd3200: data = 8'h80;
            20'd3201: data = 8'h7F;
            20'd3202: data = 8'h7F;
            20'd3203: data = 8'h80;
            20'd3204: data = 8'h80;
            20'd3205: data = 8'h80;
            20'd3206: data = 8'h7F;
            20'd3207: data = 8'h7F;
            20'd3208: data = 8'h80;
            20'd3209: data = 8'h80;
            20'd3210: data = 8'h7F;
            20'd3211: data = 8'h7F;
            20'd3212: data = 8'h80;
            20'd3213: data = 8'h7F;
            20'd3214: data = 8'h80;
            20'd3215: data = 8'h80;
            20'd3216: data = 8'h7F;
            20'd3217: data = 8'h80;
            20'd3218: data = 8'h7F;
            20'd3219: data = 8'h80;
            20'd3220: data = 8'h7F;
            20'd3221: data = 8'h80;
            20'd3222: data = 8'h7F;
            20'd3223: data = 8'h80;
            20'd3224: data = 8'h80;
            20'd3225: data = 8'h80;
            20'd3226: data = 8'h7F;
            20'd3227: data = 8'h80;
            20'd3228: data = 8'h80;
            20'd3229: data = 8'h80;
            20'd3230: data = 8'h7F;
            20'd3231: data = 8'h80;
            20'd3232: data = 8'h7F;
            20'd3233: data = 8'h7F;
            20'd3234: data = 8'h80;
            20'd3235: data = 8'h80;
            20'd3236: data = 8'h7F;
            20'd3237: data = 8'h7F;
            20'd3238: data = 8'h7F;
            20'd3239: data = 8'h80;
            20'd3240: data = 8'h7F;
            20'd3241: data = 8'h7F;
            20'd3242: data = 8'h80;
            20'd3243: data = 8'h7F;
            20'd3244: data = 8'h7F;
            20'd3245: data = 8'h7F;
            20'd3246: data = 8'h80;
            20'd3247: data = 8'h80;
            20'd3248: data = 8'h7F;
            20'd3249: data = 8'h7F;
            20'd3250: data = 8'h80;
            20'd3251: data = 8'h80;
            20'd3252: data = 8'h7F;
            20'd3253: data = 8'h80;
            20'd3254: data = 8'h7F;
            20'd3255: data = 8'h7F;
            20'd3256: data = 8'h7F;
            20'd3257: data = 8'h7F;
            20'd3258: data = 8'h7F;
            20'd3259: data = 8'h80;
            20'd3260: data = 8'h80;
            20'd3261: data = 8'h7F;
            20'd3262: data = 8'h7F;
            20'd3263: data = 8'h7F;
            20'd3264: data = 8'h80;
            20'd3265: data = 8'h7F;
            20'd3266: data = 8'h7F;
            20'd3267: data = 8'h80;
            20'd3268: data = 8'h80;
            20'd3269: data = 8'h80;
            20'd3270: data = 8'h7F;
            20'd3271: data = 8'h7F;
            20'd3272: data = 8'h7F;
            20'd3273: data = 8'h80;
            20'd3274: data = 8'h7F;
            20'd3275: data = 8'h80;
            20'd3276: data = 8'h80;
            20'd3277: data = 8'h7F;
            20'd3278: data = 8'h7F;
            20'd3279: data = 8'h7F;
            20'd3280: data = 8'h7F;
            20'd3281: data = 8'h7F;
            20'd3282: data = 8'h80;
            20'd3283: data = 8'h7F;
            20'd3284: data = 8'h80;
            20'd3285: data = 8'h80;
            20'd3286: data = 8'h80;
            20'd3287: data = 8'h7F;
            20'd3288: data = 8'h7F;
            20'd3289: data = 8'h80;
            20'd3290: data = 8'h80;
            20'd3291: data = 8'h80;
            20'd3292: data = 8'h80;
            20'd3293: data = 8'h80;
            20'd3294: data = 8'h7F;
            20'd3295: data = 8'h80;
            20'd3296: data = 8'h80;
            20'd3297: data = 8'h80;
            20'd3298: data = 8'h80;
            20'd3299: data = 8'h80;
            20'd3300: data = 8'h80;
            20'd3301: data = 8'h7F;
            20'd3302: data = 8'h80;
            20'd3303: data = 8'h80;
            20'd3304: data = 8'h80;
            20'd3305: data = 8'h80;
            20'd3306: data = 8'h80;
            20'd3307: data = 8'h80;
            20'd3308: data = 8'h80;
            20'd3309: data = 8'h80;
            20'd3310: data = 8'h7F;
            20'd3311: data = 8'h80;
            20'd3312: data = 8'h7F;
            20'd3313: data = 8'h80;
            20'd3314: data = 8'h80;
            20'd3315: data = 8'h7F;
            20'd3316: data = 8'h80;
            20'd3317: data = 8'h80;
            20'd3318: data = 8'h80;
            20'd3319: data = 8'h80;
            20'd3320: data = 8'h80;
            20'd3321: data = 8'h80;
            20'd3322: data = 8'h7F;
            20'd3323: data = 8'h80;
            20'd3324: data = 8'h80;
            20'd3325: data = 8'h80;
            20'd3326: data = 8'h80;
            20'd3327: data = 8'h80;
            20'd3328: data = 8'h80;
            20'd3329: data = 8'h80;
            20'd3330: data = 8'h80;
            20'd3331: data = 8'h80;
            20'd3332: data = 8'h7F;
            20'd3333: data = 8'h7F;
            20'd3334: data = 8'h80;
            20'd3335: data = 8'h80;
            20'd3336: data = 8'h80;
            20'd3337: data = 8'h80;
            20'd3338: data = 8'h80;
            20'd3339: data = 8'h80;
            20'd3340: data = 8'h80;
            20'd3341: data = 8'h80;
            20'd3342: data = 8'h80;
            20'd3343: data = 8'h80;
            20'd3344: data = 8'h80;
            20'd3345: data = 8'h80;
            20'd3346: data = 8'h80;
            20'd3347: data = 8'h80;
            20'd3348: data = 8'h80;
            20'd3349: data = 8'h7F;
            20'd3350: data = 8'h80;
            20'd3351: data = 8'h80;
            20'd3352: data = 8'h80;
            20'd3353: data = 8'h7F;
            20'd3354: data = 8'h80;
            20'd3355: data = 8'h80;
            20'd3356: data = 8'h80;
            20'd3357: data = 8'h7F;
            20'd3358: data = 8'h80;
            20'd3359: data = 8'h80;
            20'd3360: data = 8'h7F;
            20'd3361: data = 8'h7F;
            20'd3362: data = 8'h80;
            20'd3363: data = 8'h80;
            20'd3364: data = 8'h80;
            20'd3365: data = 8'h80;
            20'd3366: data = 8'h80;
            20'd3367: data = 8'h7F;
            20'd3368: data = 8'h80;
            20'd3369: data = 8'h80;
            20'd3370: data = 8'h7F;
            20'd3371: data = 8'h80;
            20'd3372: data = 8'h80;
            20'd3373: data = 8'h80;
            20'd3374: data = 8'h7F;
            20'd3375: data = 8'h80;
            20'd3376: data = 8'h80;
            20'd3377: data = 8'h7F;
            20'd3378: data = 8'h80;
            20'd3379: data = 8'h80;
            20'd3380: data = 8'h80;
            20'd3381: data = 8'h80;
            20'd3382: data = 8'h80;
            20'd3383: data = 8'h80;
            20'd3384: data = 8'h7F;
            20'd3385: data = 8'h80;
            20'd3386: data = 8'h7F;
            20'd3387: data = 8'h7F;
            20'd3388: data = 8'h7F;
            20'd3389: data = 8'h7F;
            20'd3390: data = 8'h80;
            20'd3391: data = 8'h80;
            20'd3392: data = 8'h80;
            20'd3393: data = 8'h80;
            20'd3394: data = 8'h80;
            20'd3395: data = 8'h7F;
            20'd3396: data = 8'h80;
            20'd3397: data = 8'h80;
            20'd3398: data = 8'h80;
            20'd3399: data = 8'h7F;
            20'd3400: data = 8'h80;
            20'd3401: data = 8'h80;
            20'd3402: data = 8'h7F;
            20'd3403: data = 8'h7F;
            20'd3404: data = 8'h7F;
            20'd3405: data = 8'h80;
            20'd3406: data = 8'h80;
            20'd3407: data = 8'h80;
            20'd3408: data = 8'h7F;
            20'd3409: data = 8'h80;
            20'd3410: data = 8'h7F;
            20'd3411: data = 8'h80;
            20'd3412: data = 8'h80;
            20'd3413: data = 8'h80;
            20'd3414: data = 8'h80;
            20'd3415: data = 8'h80;
            20'd3416: data = 8'h7F;
            20'd3417: data = 8'h7F;
            20'd3418: data = 8'h7F;
            20'd3419: data = 8'h7F;
            20'd3420: data = 8'h80;
            20'd3421: data = 8'h80;
            20'd3422: data = 8'h80;
            20'd3423: data = 8'h80;
            20'd3424: data = 8'h80;
            20'd3425: data = 8'h7F;
            20'd3426: data = 8'h7F;
            20'd3427: data = 8'h80;
            20'd3428: data = 8'h7F;
            20'd3429: data = 8'h80;
            20'd3430: data = 8'h7F;
            20'd3431: data = 8'h80;
            20'd3432: data = 8'h80;
            20'd3433: data = 8'h80;
            20'd3434: data = 8'h7F;
            20'd3435: data = 8'h80;
            20'd3436: data = 8'h80;
            20'd3437: data = 8'h80;
            20'd3438: data = 8'h80;
            20'd3439: data = 8'h80;
            20'd3440: data = 8'h80;
            20'd3441: data = 8'h7F;
            20'd3442: data = 8'h80;
            20'd3443: data = 8'h7F;
            20'd3444: data = 8'h80;
            20'd3445: data = 8'h80;
            20'd3446: data = 8'h80;
            20'd3447: data = 8'h80;
            20'd3448: data = 8'h80;
            20'd3449: data = 8'h80;
            20'd3450: data = 8'h80;
            20'd3451: data = 8'h80;
            20'd3452: data = 8'h80;
            20'd3453: data = 8'h80;
            20'd3454: data = 8'h80;
            20'd3455: data = 8'h80;
            20'd3456: data = 8'h7F;
            20'd3457: data = 8'h7F;
            20'd3458: data = 8'h80;
            20'd3459: data = 8'h80;
            20'd3460: data = 8'h80;
            20'd3461: data = 8'h80;
            20'd3462: data = 8'h80;
            20'd3463: data = 8'h80;
            20'd3464: data = 8'h7F;
            20'd3465: data = 8'h80;
            20'd3466: data = 8'h80;
            20'd3467: data = 8'h7F;
            20'd3468: data = 8'h7F;
            20'd3469: data = 8'h7F;
            20'd3470: data = 8'h80;
            20'd3471: data = 8'h80;
            20'd3472: data = 8'h80;
            20'd3473: data = 8'h80;
            20'd3474: data = 8'h7F;
            20'd3475: data = 8'h80;
            20'd3476: data = 8'h7F;
            20'd3477: data = 8'h7F;
            20'd3478: data = 8'h80;
            20'd3479: data = 8'h80;
            20'd3480: data = 8'h80;
            20'd3481: data = 8'h80;
            20'd3482: data = 8'h80;
            20'd3483: data = 8'h80;
            20'd3484: data = 8'h80;
            20'd3485: data = 8'h7F;
            20'd3486: data = 8'h80;
            20'd3487: data = 8'h80;
            20'd3488: data = 8'h80;
            20'd3489: data = 8'h80;
            20'd3490: data = 8'h80;
            20'd3491: data = 8'h80;
            20'd3492: data = 8'h80;
            20'd3493: data = 8'h7F;
            20'd3494: data = 8'h80;
            20'd3495: data = 8'h80;
            20'd3496: data = 8'h80;
            20'd3497: data = 8'h80;
            20'd3498: data = 8'h80;
            20'd3499: data = 8'h80;
            20'd3500: data = 8'h80;
            20'd3501: data = 8'h7F;
            20'd3502: data = 8'h7F;
            20'd3503: data = 8'h7F;
            20'd3504: data = 8'h80;
            20'd3505: data = 8'h80;
            20'd3506: data = 8'h80;
            20'd3507: data = 8'h80;
            20'd3508: data = 8'h7F;
            20'd3509: data = 8'h7F;
            20'd3510: data = 8'h80;
            20'd3511: data = 8'h80;
            20'd3512: data = 8'h80;
            20'd3513: data = 8'h80;
            20'd3514: data = 8'h80;
            20'd3515: data = 8'h80;
            20'd3516: data = 8'h80;
            20'd3517: data = 8'h80;
            20'd3518: data = 8'h7F;
            20'd3519: data = 8'h7F;
            20'd3520: data = 8'h80;
            20'd3521: data = 8'h7F;
            20'd3522: data = 8'h7F;
            20'd3523: data = 8'h80;
            20'd3524: data = 8'h80;
            20'd3525: data = 8'h80;
            20'd3526: data = 8'h80;
            20'd3527: data = 8'h7F;
            20'd3528: data = 8'h80;
            20'd3529: data = 8'h80;
            20'd3530: data = 8'h80;
            20'd3531: data = 8'h7F;
            20'd3532: data = 8'h80;
            20'd3533: data = 8'h80;
            20'd3534: data = 8'h80;
            20'd3535: data = 8'h80;
            20'd3536: data = 8'h7F;
            20'd3537: data = 8'h80;
            20'd3538: data = 8'h80;
            20'd3539: data = 8'h80;
            20'd3540: data = 8'h80;
            20'd3541: data = 8'h80;
            20'd3542: data = 8'h7F;
            20'd3543: data = 8'h7F;
            20'd3544: data = 8'h80;
            20'd3545: data = 8'h80;
            20'd3546: data = 8'h80;
            20'd3547: data = 8'h80;
            20'd3548: data = 8'h7F;
            20'd3549: data = 8'h80;
            20'd3550: data = 8'h80;
            20'd3551: data = 8'h80;
            20'd3552: data = 8'h7F;
            20'd3553: data = 8'h7F;
            20'd3554: data = 8'h80;
            20'd3555: data = 8'h80;
            20'd3556: data = 8'h80;
            20'd3557: data = 8'h80;
            20'd3558: data = 8'h80;
            20'd3559: data = 8'h80;
            20'd3560: data = 8'h80;
            20'd3561: data = 8'h80;
            20'd3562: data = 8'h7F;
            20'd3563: data = 8'h80;
            20'd3564: data = 8'h80;
            20'd3565: data = 8'h80;
            20'd3566: data = 8'h80;
            20'd3567: data = 8'h7F;
            20'd3568: data = 8'h7F;
            20'd3569: data = 8'h80;
            20'd3570: data = 8'h80;
            20'd3571: data = 8'h80;
            20'd3572: data = 8'h7F;
            20'd3573: data = 8'h80;
            20'd3574: data = 8'h7F;
            20'd3575: data = 8'h7F;
            20'd3576: data = 8'h7F;
            20'd3577: data = 8'h80;
            20'd3578: data = 8'h80;
            20'd3579: data = 8'h80;
            20'd3580: data = 8'h80;
            20'd3581: data = 8'h80;
            20'd3582: data = 8'h80;
            20'd3583: data = 8'h80;
            20'd3584: data = 8'h80;
            20'd3585: data = 8'h80;
            20'd3586: data = 8'h80;
            20'd3587: data = 8'h80;
            20'd3588: data = 8'h80;
            20'd3589: data = 8'h80;
            20'd3590: data = 8'h80;
            20'd3591: data = 8'h7F;
            20'd3592: data = 8'h7F;
            20'd3593: data = 8'h80;
            20'd3594: data = 8'h7F;
            20'd3595: data = 8'h80;
            20'd3596: data = 8'h80;
            20'd3597: data = 8'h80;
            20'd3598: data = 8'h80;
            20'd3599: data = 8'h7F;
            20'd3600: data = 8'h80;
            20'd3601: data = 8'h80;
            20'd3602: data = 8'h80;
            20'd3603: data = 8'h80;
            20'd3604: data = 8'h7F;
            20'd3605: data = 8'h80;
            20'd3606: data = 8'h80;
            20'd3607: data = 8'h80;
            20'd3608: data = 8'h7F;
            20'd3609: data = 8'h80;
            20'd3610: data = 8'h80;
            20'd3611: data = 8'h80;
            20'd3612: data = 8'h80;
            20'd3613: data = 8'h7F;
            20'd3614: data = 8'h7F;
            20'd3615: data = 8'h7F;
            20'd3616: data = 8'h80;
            20'd3617: data = 8'h7F;
            20'd3618: data = 8'h7F;
            20'd3619: data = 8'h80;
            20'd3620: data = 8'h80;
            20'd3621: data = 8'h80;
            20'd3622: data = 8'h7F;
            20'd3623: data = 8'h80;
            20'd3624: data = 8'h80;
            20'd3625: data = 8'h80;
            20'd3626: data = 8'h80;
            20'd3627: data = 8'h80;
            20'd3628: data = 8'h80;
            20'd3629: data = 8'h80;
            20'd3630: data = 8'h80;
            20'd3631: data = 8'h80;
            20'd3632: data = 8'h80;
            20'd3633: data = 8'h80;
            20'd3634: data = 8'h80;
            20'd3635: data = 8'h7F;
            20'd3636: data = 8'h80;
            20'd3637: data = 8'h80;
            20'd3638: data = 8'h7F;
            20'd3639: data = 8'h80;
            20'd3640: data = 8'h7F;
            20'd3641: data = 8'h80;
            20'd3642: data = 8'h80;
            20'd3643: data = 8'h80;
            20'd3644: data = 8'h7F;
            20'd3645: data = 8'h80;
            20'd3646: data = 8'h7F;
            20'd3647: data = 8'h80;
            20'd3648: data = 8'h80;
            20'd3649: data = 8'h80;
            20'd3650: data = 8'h80;
            20'd3651: data = 8'h80;
            20'd3652: data = 8'h7F;
            20'd3653: data = 8'h7F;
            20'd3654: data = 8'h80;
            20'd3655: data = 8'h80;
            20'd3656: data = 8'h80;
            20'd3657: data = 8'h80;
            20'd3658: data = 8'h80;
            20'd3659: data = 8'h80;
            20'd3660: data = 8'h7F;
            20'd3661: data = 8'h80;
            20'd3662: data = 8'h80;
            20'd3663: data = 8'h7F;
            20'd3664: data = 8'h80;
            20'd3665: data = 8'h7F;
            20'd3666: data = 8'h7F;
            20'd3667: data = 8'h80;
            20'd3668: data = 8'h80;
            20'd3669: data = 8'h80;
            20'd3670: data = 8'h80;
            20'd3671: data = 8'h80;
            20'd3672: data = 8'h80;
            20'd3673: data = 8'h80;
            20'd3674: data = 8'h80;
            20'd3675: data = 8'h7F;
            20'd3676: data = 8'h7F;
            20'd3677: data = 8'h80;
            20'd3678: data = 8'h7F;
            20'd3679: data = 8'h80;
            20'd3680: data = 8'h7F;
            20'd3681: data = 8'h80;
            20'd3682: data = 8'h80;
            20'd3683: data = 8'h80;
            20'd3684: data = 8'h7F;
            20'd3685: data = 8'h7F;
            20'd3686: data = 8'h80;
            20'd3687: data = 8'h7F;
            20'd3688: data = 8'h7F;
            20'd3689: data = 8'h7F;
            20'd3690: data = 8'h80;
            20'd3691: data = 8'h7F;
            20'd3692: data = 8'h80;
            20'd3693: data = 8'h80;
            20'd3694: data = 8'h7F;
            20'd3695: data = 8'h7F;
            20'd3696: data = 8'h7F;
            20'd3697: data = 8'h80;
            20'd3698: data = 8'h80;
            20'd3699: data = 8'h7F;
            20'd3700: data = 8'h80;
            20'd3701: data = 8'h7F;
            20'd3702: data = 8'h80;
            20'd3703: data = 8'h80;
            20'd3704: data = 8'h80;
            20'd3705: data = 8'h7F;
            20'd3706: data = 8'h80;
            20'd3707: data = 8'h80;
            20'd3708: data = 8'h80;
            20'd3709: data = 8'h7F;
            20'd3710: data = 8'h80;
            20'd3711: data = 8'h80;
            20'd3712: data = 8'h80;
            20'd3713: data = 8'h7F;
            20'd3714: data = 8'h80;
            20'd3715: data = 8'h80;
            20'd3716: data = 8'h80;
            20'd3717: data = 8'h80;
            20'd3718: data = 8'h80;
            20'd3719: data = 8'h7F;
            20'd3720: data = 8'h80;
            20'd3721: data = 8'h80;
            20'd3722: data = 8'h80;
            20'd3723: data = 8'h80;
            20'd3724: data = 8'h80;
            20'd3725: data = 8'h7F;
            20'd3726: data = 8'h80;
            20'd3727: data = 8'h80;
            20'd3728: data = 8'h7F;
            20'd3729: data = 8'h80;
            20'd3730: data = 8'h80;
            20'd3731: data = 8'h80;
            20'd3732: data = 8'h80;
            20'd3733: data = 8'h7F;
            20'd3734: data = 8'h80;
            20'd3735: data = 8'h80;
            20'd3736: data = 8'h7F;
            20'd3737: data = 8'h80;
            20'd3738: data = 8'h80;
            20'd3739: data = 8'h80;
            20'd3740: data = 8'h80;
            20'd3741: data = 8'h7F;
            20'd3742: data = 8'h7F;
            20'd3743: data = 8'h80;
            20'd3744: data = 8'h80;
            20'd3745: data = 8'h80;
            20'd3746: data = 8'h80;
            20'd3747: data = 8'h80;
            20'd3748: data = 8'h7F;
            20'd3749: data = 8'h7F;
            20'd3750: data = 8'h80;
            20'd3751: data = 8'h80;
            20'd3752: data = 8'h7F;
            20'd3753: data = 8'h80;
            20'd3754: data = 8'h7F;
            20'd3755: data = 8'h7F;
            20'd3756: data = 8'h80;
            20'd3757: data = 8'h80;
            20'd3758: data = 8'h80;
            20'd3759: data = 8'h7F;
            20'd3760: data = 8'h80;
            20'd3761: data = 8'h80;
            20'd3762: data = 8'h80;
            20'd3763: data = 8'h7F;
            20'd3764: data = 8'h7F;
            20'd3765: data = 8'h80;
            20'd3766: data = 8'h80;
            20'd3767: data = 8'h80;
            20'd3768: data = 8'h80;
            20'd3769: data = 8'h7F;
            20'd3770: data = 8'h80;
            20'd3771: data = 8'h80;
            20'd3772: data = 8'h80;
            20'd3773: data = 8'h7F;
            20'd3774: data = 8'h80;
            20'd3775: data = 8'h80;
            20'd3776: data = 8'h80;
            20'd3777: data = 8'h80;
            20'd3778: data = 8'h80;
            20'd3779: data = 8'h80;
            20'd3780: data = 8'h7F;
            20'd3781: data = 8'h80;
            20'd3782: data = 8'h80;
            20'd3783: data = 8'h7F;
            20'd3784: data = 8'h80;
            20'd3785: data = 8'h80;
            20'd3786: data = 8'h7F;
            20'd3787: data = 8'h80;
            20'd3788: data = 8'h80;
            20'd3789: data = 8'h7F;
            20'd3790: data = 8'h80;
            20'd3791: data = 8'h80;
            20'd3792: data = 8'h7F;
            20'd3793: data = 8'h80;
            20'd3794: data = 8'h80;
            20'd3795: data = 8'h80;
            20'd3796: data = 8'h80;
            20'd3797: data = 8'h7F;
            20'd3798: data = 8'h7F;
            20'd3799: data = 8'h7F;
            20'd3800: data = 8'h80;
            20'd3801: data = 8'h80;
            20'd3802: data = 8'h7F;
            20'd3803: data = 8'h80;
            20'd3804: data = 8'h80;
            20'd3805: data = 8'h80;
            20'd3806: data = 8'h80;
            20'd3807: data = 8'h7F;
            20'd3808: data = 8'h80;
            20'd3809: data = 8'h80;
            20'd3810: data = 8'h7F;
            20'd3811: data = 8'h80;
            20'd3812: data = 8'h7F;
            20'd3813: data = 8'h80;
            20'd3814: data = 8'h80;
            20'd3815: data = 8'h80;
            20'd3816: data = 8'h80;
            20'd3817: data = 8'h80;
            20'd3818: data = 8'h80;
            20'd3819: data = 8'h7F;
            20'd3820: data = 8'h80;
            20'd3821: data = 8'h80;
            20'd3822: data = 8'h7F;
            20'd3823: data = 8'h7F;
            20'd3824: data = 8'h80;
            20'd3825: data = 8'h80;
            20'd3826: data = 8'h80;
            20'd3827: data = 8'h80;
            20'd3828: data = 8'h7F;
            20'd3829: data = 8'h7F;
            20'd3830: data = 8'h80;
            20'd3831: data = 8'h7F;
            20'd3832: data = 8'h80;
            20'd3833: data = 8'h7F;
            20'd3834: data = 8'h7F;
            20'd3835: data = 8'h80;
            20'd3836: data = 8'h7F;
            20'd3837: data = 8'h7F;
            20'd3838: data = 8'h80;
            20'd3839: data = 8'h7F;
            20'd3840: data = 8'h7F;
            20'd3841: data = 8'h80;
            20'd3842: data = 8'h80;
            20'd3843: data = 8'h80;
            20'd3844: data = 8'h80;
            20'd3845: data = 8'h7F;
            20'd3846: data = 8'h80;
            20'd3847: data = 8'h80;
            20'd3848: data = 8'h80;
            20'd3849: data = 8'h80;
            20'd3850: data = 8'h80;
            20'd3851: data = 8'h7F;
            20'd3852: data = 8'h80;
            20'd3853: data = 8'h7F;
            20'd3854: data = 8'h7F;
            20'd3855: data = 8'h80;
            20'd3856: data = 8'h80;
            20'd3857: data = 8'h80;
            20'd3858: data = 8'h7F;
            20'd3859: data = 8'h80;
            20'd3860: data = 8'h80;
            20'd3861: data = 8'h7F;
            20'd3862: data = 8'h7F;
            20'd3863: data = 8'h80;
            20'd3864: data = 8'h80;
            20'd3865: data = 8'h7F;
            20'd3866: data = 8'h80;
            20'd3867: data = 8'h80;
            20'd3868: data = 8'h80;
            20'd3869: data = 8'h80;
            20'd3870: data = 8'h80;
            20'd3871: data = 8'h80;
            20'd3872: data = 8'h7F;
            20'd3873: data = 8'h80;
            20'd3874: data = 8'h7F;
            20'd3875: data = 8'h80;
            20'd3876: data = 8'h7F;
            20'd3877: data = 8'h7F;
            20'd3878: data = 8'h80;
            20'd3879: data = 8'h7F;
            20'd3880: data = 8'h80;
            20'd3881: data = 8'h80;
            20'd3882: data = 8'h80;
            20'd3883: data = 8'h7F;
            20'd3884: data = 8'h80;
            20'd3885: data = 8'h80;
            20'd3886: data = 8'h80;
            20'd3887: data = 8'h7F;
            20'd3888: data = 8'h80;
            20'd3889: data = 8'h80;
            20'd3890: data = 8'h7F;
            20'd3891: data = 8'h7F;
            20'd3892: data = 8'h80;
            20'd3893: data = 8'h7F;
            20'd3894: data = 8'h80;
            20'd3895: data = 8'h80;
            20'd3896: data = 8'h80;
            20'd3897: data = 8'h80;
            20'd3898: data = 8'h7F;
            20'd3899: data = 8'h80;
            20'd3900: data = 8'h80;
            20'd3901: data = 8'h80;
            20'd3902: data = 8'h80;
            20'd3903: data = 8'h80;
            20'd3904: data = 8'h7F;
            20'd3905: data = 8'h7F;
            20'd3906: data = 8'h80;
            20'd3907: data = 8'h80;
            20'd3908: data = 8'h80;
            20'd3909: data = 8'h7F;
            20'd3910: data = 8'h80;
            20'd3911: data = 8'h80;
            20'd3912: data = 8'h7F;
            20'd3913: data = 8'h80;
            20'd3914: data = 8'h80;
            20'd3915: data = 8'h7F;
            20'd3916: data = 8'h80;
            20'd3917: data = 8'h80;
            20'd3918: data = 8'h7F;
            20'd3919: data = 8'h80;
            20'd3920: data = 8'h7F;
            20'd3921: data = 8'h7F;
            20'd3922: data = 8'h7F;
            20'd3923: data = 8'h7F;
            20'd3924: data = 8'h80;
            20'd3925: data = 8'h7F;
            20'd3926: data = 8'h80;
            20'd3927: data = 8'h80;
            20'd3928: data = 8'h80;
            20'd3929: data = 8'h80;
            20'd3930: data = 8'h7F;
            20'd3931: data = 8'h80;
            20'd3932: data = 8'h80;
            20'd3933: data = 8'h80;
            20'd3934: data = 8'h80;
            20'd3935: data = 8'h80;
            20'd3936: data = 8'h80;
            20'd3937: data = 8'h7F;
            20'd3938: data = 8'h80;
            20'd3939: data = 8'h7F;
            20'd3940: data = 8'h80;
            20'd3941: data = 8'h7F;
            20'd3942: data = 8'h80;
            20'd3943: data = 8'h80;
            20'd3944: data = 8'h7F;
            20'd3945: data = 8'h80;
            20'd3946: data = 8'h80;
            20'd3947: data = 8'h80;
            20'd3948: data = 8'h7F;
            20'd3949: data = 8'h7F;
            20'd3950: data = 8'h7F;
            20'd3951: data = 8'h80;
            20'd3952: data = 8'h80;
            20'd3953: data = 8'h80;
            20'd3954: data = 8'h80;
            20'd3955: data = 8'h7F;
            20'd3956: data = 8'h7F;
            20'd3957: data = 8'h80;
            20'd3958: data = 8'h80;
            20'd3959: data = 8'h7F;
            20'd3960: data = 8'h80;
            20'd3961: data = 8'h80;
            20'd3962: data = 8'h80;
            20'd3963: data = 8'h80;
            20'd3964: data = 8'h80;
            20'd3965: data = 8'h7F;
            20'd3966: data = 8'h80;
            20'd3967: data = 8'h80;
            20'd3968: data = 8'h80;
            20'd3969: data = 8'h7F;
            20'd3970: data = 8'h80;
            20'd3971: data = 8'h7F;
            20'd3972: data = 8'h80;
            20'd3973: data = 8'h80;
            20'd3974: data = 8'h80;
            20'd3975: data = 8'h7F;
            20'd3976: data = 8'h80;
            20'd3977: data = 8'h80;
            20'd3978: data = 8'h80;
            20'd3979: data = 8'h80;
            20'd3980: data = 8'h7F;
            20'd3981: data = 8'h80;
            20'd3982: data = 8'h7F;
            20'd3983: data = 8'h80;
            20'd3984: data = 8'h80;
            20'd3985: data = 8'h80;
            20'd3986: data = 8'h7F;
            20'd3987: data = 8'h80;
            20'd3988: data = 8'h80;
            20'd3989: data = 8'h80;
            20'd3990: data = 8'h80;
            20'd3991: data = 8'h7F;
            20'd3992: data = 8'h7F;
            20'd3993: data = 8'h80;
            20'd3994: data = 8'h80;
            20'd3995: data = 8'h80;
            20'd3996: data = 8'h80;
            20'd3997: data = 8'h80;
            20'd3998: data = 8'h80;
            20'd3999: data = 8'h7F;
            20'd4000: data = 8'h80;
            20'd4001: data = 8'h80;
            20'd4002: data = 8'h80;
            20'd4003: data = 8'h80;
            20'd4004: data = 8'h7F;
            20'd4005: data = 8'h7F;
            20'd4006: data = 8'h7F;
            20'd4007: data = 8'h80;
            20'd4008: data = 8'h80;
            20'd4009: data = 8'h7F;
            20'd4010: data = 8'h80;
            20'd4011: data = 8'h80;
            20'd4012: data = 8'h7F;
            20'd4013: data = 8'h80;
            20'd4014: data = 8'h80;
            20'd4015: data = 8'h7F;
            20'd4016: data = 8'h80;
            20'd4017: data = 8'h80;
            20'd4018: data = 8'h7F;
            20'd4019: data = 8'h80;
            20'd4020: data = 8'h7F;
            20'd4021: data = 8'h80;
            20'd4022: data = 8'h80;
            20'd4023: data = 8'h7F;
            20'd4024: data = 8'h80;
            20'd4025: data = 8'h80;
            20'd4026: data = 8'h80;
            20'd4027: data = 8'h80;
            20'd4028: data = 8'h80;
            20'd4029: data = 8'h80;
            20'd4030: data = 8'h80;
            20'd4031: data = 8'h80;
            20'd4032: data = 8'h80;
            20'd4033: data = 8'h7F;
            20'd4034: data = 8'h80;
            20'd4035: data = 8'h80;
            20'd4036: data = 8'h7F;
            20'd4037: data = 8'h80;
            20'd4038: data = 8'h80;
            20'd4039: data = 8'h80;
            20'd4040: data = 8'h80;
            20'd4041: data = 8'h80;
            20'd4042: data = 8'h7F;
            20'd4043: data = 8'h80;
            20'd4044: data = 8'h80;
            20'd4045: data = 8'h80;
            20'd4046: data = 8'h80;
            20'd4047: data = 8'h7F;
            20'd4048: data = 8'h80;
            20'd4049: data = 8'h80;
            20'd4050: data = 8'h7F;
            20'd4051: data = 8'h80;
            20'd4052: data = 8'h7F;
            20'd4053: data = 8'h80;
            20'd4054: data = 8'h80;
            20'd4055: data = 8'h80;
            20'd4056: data = 8'h80;
            20'd4057: data = 8'h80;
            20'd4058: data = 8'h80;
            20'd4059: data = 8'h7F;
            20'd4060: data = 8'h80;
            20'd4061: data = 8'h80;
            20'd4062: data = 8'h80;
            20'd4063: data = 8'h80;
            20'd4064: data = 8'h80;
            20'd4065: data = 8'h7F;
            20'd4066: data = 8'h80;
            20'd4067: data = 8'h7F;
            20'd4068: data = 8'h80;
            20'd4069: data = 8'h80;
            20'd4070: data = 8'h80;
            20'd4071: data = 8'h7F;
            20'd4072: data = 8'h80;
            20'd4073: data = 8'h80;
            20'd4074: data = 8'h7F;
            20'd4075: data = 8'h80;
            20'd4076: data = 8'h7F;
            20'd4077: data = 8'h80;
            20'd4078: data = 8'h80;
            20'd4079: data = 8'h80;
            20'd4080: data = 8'h80;
            20'd4081: data = 8'h80;
            20'd4082: data = 8'h7F;
            20'd4083: data = 8'h80;
            20'd4084: data = 8'h80;
            20'd4085: data = 8'h80;
            20'd4086: data = 8'h80;
            20'd4087: data = 8'h7F;
            20'd4088: data = 8'h7F;
            20'd4089: data = 8'h7F;
            20'd4090: data = 8'h80;
            20'd4091: data = 8'h80;
            20'd4092: data = 8'h80;
            20'd4093: data = 8'h80;
            20'd4094: data = 8'h80;
            20'd4095: data = 8'h80;
            20'd4096: data = 8'h7F;
            20'd4097: data = 8'h80;
            20'd4098: data = 8'h80;
            20'd4099: data = 8'h80;
            20'd4100: data = 8'h7F;
            20'd4101: data = 8'h80;
            20'd4102: data = 8'h80;
            20'd4103: data = 8'h7F;
            20'd4104: data = 8'h80;
            20'd4105: data = 8'h80;
            20'd4106: data = 8'h80;
            20'd4107: data = 8'h7F;
            20'd4108: data = 8'h80;
            20'd4109: data = 8'h80;
            20'd4110: data = 8'h80;
            20'd4111: data = 8'h80;
            20'd4112: data = 8'h7F;
            20'd4113: data = 8'h7F;
            20'd4114: data = 8'h7F;
            20'd4115: data = 8'h7F;
            20'd4116: data = 8'h80;
            20'd4117: data = 8'h80;
            20'd4118: data = 8'h80;
            20'd4119: data = 8'h7F;
            20'd4120: data = 8'h80;
            20'd4121: data = 8'h80;
            20'd4122: data = 8'h80;
            20'd4123: data = 8'h80;
            20'd4124: data = 8'h7F;
            20'd4125: data = 8'h80;
            20'd4126: data = 8'h7F;
            20'd4127: data = 8'h80;
            20'd4128: data = 8'h80;
            20'd4129: data = 8'h7F;
            20'd4130: data = 8'h80;
            20'd4131: data = 8'h80;
            20'd4132: data = 8'h80;
            20'd4133: data = 8'h7F;
            20'd4134: data = 8'h80;
            20'd4135: data = 8'h7F;
            20'd4136: data = 8'h7F;
            20'd4137: data = 8'h80;
            20'd4138: data = 8'h80;
            20'd4139: data = 8'h7F;
            20'd4140: data = 8'h80;
            20'd4141: data = 8'h80;
            20'd4142: data = 8'h80;
            20'd4143: data = 8'h7F;
            20'd4144: data = 8'h80;
            20'd4145: data = 8'h7F;
            20'd4146: data = 8'h80;
            20'd4147: data = 8'h7F;
            20'd4148: data = 8'h80;
            20'd4149: data = 8'h7F;
            20'd4150: data = 8'h7F;
            20'd4151: data = 8'h80;
            20'd4152: data = 8'h80;
            20'd4153: data = 8'h7F;
            20'd4154: data = 8'h7F;
            20'd4155: data = 8'h80;
            20'd4156: data = 8'h80;
            20'd4157: data = 8'h80;
            20'd4158: data = 8'h7F;
            20'd4159: data = 8'h80;
            20'd4160: data = 8'h7F;
            20'd4161: data = 8'h80;
            20'd4162: data = 8'h80;
            20'd4163: data = 8'h7F;
            20'd4164: data = 8'h80;
            20'd4165: data = 8'h80;
            20'd4166: data = 8'h7F;
            20'd4167: data = 8'h80;
            20'd4168: data = 8'h80;
            20'd4169: data = 8'h7F;
            20'd4170: data = 8'h80;
            20'd4171: data = 8'h80;
            20'd4172: data = 8'h7F;
            20'd4173: data = 8'h80;
            20'd4174: data = 8'h80;
            20'd4175: data = 8'h7F;
            20'd4176: data = 8'h7F;
            20'd4177: data = 8'h80;
            20'd4178: data = 8'h7F;
            20'd4179: data = 8'h7F;
            20'd4180: data = 8'h7F;
            20'd4181: data = 8'h80;
            20'd4182: data = 8'h80;
            20'd4183: data = 8'h80;
            20'd4184: data = 8'h80;
            20'd4185: data = 8'h7F;
            20'd4186: data = 8'h80;
            20'd4187: data = 8'h80;
            20'd4188: data = 8'h80;
            20'd4189: data = 8'h7F;
            20'd4190: data = 8'h7F;
            20'd4191: data = 8'h80;
            20'd4192: data = 8'h80;
            20'd4193: data = 8'h80;
            20'd4194: data = 8'h80;
            20'd4195: data = 8'h80;
            20'd4196: data = 8'h80;
            20'd4197: data = 8'h7F;
            20'd4198: data = 8'h80;
            20'd4199: data = 8'h80;
            20'd4200: data = 8'h7F;
            20'd4201: data = 8'h7F;
            20'd4202: data = 8'h80;
            20'd4203: data = 8'h80;
            20'd4204: data = 8'h80;
            20'd4205: data = 8'h80;
            20'd4206: data = 8'h80;
            20'd4207: data = 8'h7F;
            20'd4208: data = 8'h7F;
            20'd4209: data = 8'h80;
            20'd4210: data = 8'h7F;
            20'd4211: data = 8'h7F;
            20'd4212: data = 8'h7F;
            20'd4213: data = 8'h7F;
            20'd4214: data = 8'h80;
            20'd4215: data = 8'h80;
            20'd4216: data = 8'h7F;
            20'd4217: data = 8'h7F;
            20'd4218: data = 8'h7F;
            20'd4219: data = 8'h7F;
            20'd4220: data = 8'h80;
            20'd4221: data = 8'h80;
            20'd4222: data = 8'h7F;
            20'd4223: data = 8'h80;
            20'd4224: data = 8'h7F;
            20'd4225: data = 8'h80;
            20'd4226: data = 8'h80;
            20'd4227: data = 8'h80;
            20'd4228: data = 8'h80;
            20'd4229: data = 8'h7F;
            20'd4230: data = 8'h80;
            20'd4231: data = 8'h80;
            20'd4232: data = 8'h80;
            20'd4233: data = 8'h80;
            20'd4234: data = 8'h80;
            20'd4235: data = 8'h7F;
            20'd4236: data = 8'h80;
            20'd4237: data = 8'h7F;
            20'd4238: data = 8'h80;
            20'd4239: data = 8'h80;
            20'd4240: data = 8'h80;
            20'd4241: data = 8'h7F;
            20'd4242: data = 8'h7F;
            20'd4243: data = 8'h80;
            20'd4244: data = 8'h80;
            20'd4245: data = 8'h7F;
            20'd4246: data = 8'h7F;
            20'd4247: data = 8'h7F;
            20'd4248: data = 8'h80;
            20'd4249: data = 8'h80;
            20'd4250: data = 8'h80;
            20'd4251: data = 8'h80;
            20'd4252: data = 8'h80;
            20'd4253: data = 8'h80;
            20'd4254: data = 8'h7F;
            20'd4255: data = 8'h80;
            20'd4256: data = 8'h7F;
            20'd4257: data = 8'h80;
            20'd4258: data = 8'h80;
            20'd4259: data = 8'h7F;
            20'd4260: data = 8'h80;
            20'd4261: data = 8'h7F;
            20'd4262: data = 8'h80;
            20'd4263: data = 8'h80;
            20'd4264: data = 8'h7F;
            20'd4265: data = 8'h80;
            20'd4266: data = 8'h7F;
            20'd4267: data = 8'h80;
            20'd4268: data = 8'h7F;
            20'd4269: data = 8'h80;
            20'd4270: data = 8'h80;
            20'd4271: data = 8'h80;
            20'd4272: data = 8'h80;
            20'd4273: data = 8'h80;
            20'd4274: data = 8'h80;
            20'd4275: data = 8'h80;
            20'd4276: data = 8'h80;
            20'd4277: data = 8'h80;
            20'd4278: data = 8'h80;
            20'd4279: data = 8'h80;
            20'd4280: data = 8'h7F;
            20'd4281: data = 8'h80;
            20'd4282: data = 8'h7F;
            20'd4283: data = 8'h80;
            20'd4284: data = 8'h7F;
            20'd4285: data = 8'h7F;
            20'd4286: data = 8'h80;
            20'd4287: data = 8'h80;
            20'd4288: data = 8'h80;
            20'd4289: data = 8'h7F;
            20'd4290: data = 8'h7F;
            20'd4291: data = 8'h80;
            20'd4292: data = 8'h80;
            20'd4293: data = 8'h7F;
            20'd4294: data = 8'h7F;
            20'd4295: data = 8'h7F;
            20'd4296: data = 8'h7F;
            20'd4297: data = 8'h80;
            20'd4298: data = 8'h80;
            20'd4299: data = 8'h80;
            20'd4300: data = 8'h7F;
            20'd4301: data = 8'h80;
            20'd4302: data = 8'h7F;
            20'd4303: data = 8'h80;
            20'd4304: data = 8'h7F;
            20'd4305: data = 8'h80;
            20'd4306: data = 8'h80;
            20'd4307: data = 8'h80;
            20'd4308: data = 8'h80;
            20'd4309: data = 8'h7F;
            20'd4310: data = 8'h80;
            20'd4311: data = 8'h80;
            20'd4312: data = 8'h7F;
            20'd4313: data = 8'h80;
            20'd4314: data = 8'h7F;
            20'd4315: data = 8'h7F;
            20'd4316: data = 8'h80;
            20'd4317: data = 8'h80;
            20'd4318: data = 8'h80;
            20'd4319: data = 8'h80;
            20'd4320: data = 8'h80;
            20'd4321: data = 8'h80;
            20'd4322: data = 8'h7F;
            20'd4323: data = 8'h80;
            20'd4324: data = 8'h7F;
            20'd4325: data = 8'h80;
            20'd4326: data = 8'h80;
            20'd4327: data = 8'h7F;
            20'd4328: data = 8'h80;
            20'd4329: data = 8'h80;
            20'd4330: data = 8'h80;
            20'd4331: data = 8'h80;
            20'd4332: data = 8'h80;
            20'd4333: data = 8'h80;
            20'd4334: data = 8'h80;
            20'd4335: data = 8'h80;
            20'd4336: data = 8'h80;
            20'd4337: data = 8'h80;
            20'd4338: data = 8'h7F;
            20'd4339: data = 8'h7F;
            20'd4340: data = 8'h80;
            20'd4341: data = 8'h80;
            20'd4342: data = 8'h80;
            20'd4343: data = 8'h7F;
            20'd4344: data = 8'h80;
            20'd4345: data = 8'h80;
            20'd4346: data = 8'h80;
            20'd4347: data = 8'h80;
            20'd4348: data = 8'h80;
            20'd4349: data = 8'h80;
            20'd4350: data = 8'h80;
            20'd4351: data = 8'h7F;
            20'd4352: data = 8'h80;
            20'd4353: data = 8'h80;
            20'd4354: data = 8'h7F;
            20'd4355: data = 8'h7F;
            20'd4356: data = 8'h80;
            20'd4357: data = 8'h80;
            20'd4358: data = 8'h7F;
            20'd4359: data = 8'h80;
            20'd4360: data = 8'h80;
            20'd4361: data = 8'h7F;
            20'd4362: data = 8'h7F;
            20'd4363: data = 8'h80;
            20'd4364: data = 8'h7F;
            20'd4365: data = 8'h7F;
            20'd4366: data = 8'h80;
            20'd4367: data = 8'h7F;
            20'd4368: data = 8'h80;
            20'd4369: data = 8'h7F;
            20'd4370: data = 8'h80;
            20'd4371: data = 8'h7F;
            20'd4372: data = 8'h7F;
            20'd4373: data = 8'h80;
            20'd4374: data = 8'h80;
            20'd4375: data = 8'h80;
            20'd4376: data = 8'h7F;
            20'd4377: data = 8'h80;
            20'd4378: data = 8'h7F;
            20'd4379: data = 8'h7F;
            20'd4380: data = 8'h7F;
            20'd4381: data = 8'h80;
            20'd4382: data = 8'h80;
            20'd4383: data = 8'h7F;
            20'd4384: data = 8'h7F;
            20'd4385: data = 8'h7F;
            20'd4386: data = 8'h80;
            20'd4387: data = 8'h80;
            20'd4388: data = 8'h7F;
            20'd4389: data = 8'h80;
            20'd4390: data = 8'h80;
            20'd4391: data = 8'h7F;
            20'd4392: data = 8'h80;
            20'd4393: data = 8'h80;
            20'd4394: data = 8'h7F;
            20'd4395: data = 8'h7F;
            20'd4396: data = 8'h80;
            20'd4397: data = 8'h80;
            20'd4398: data = 8'h80;
            20'd4399: data = 8'h7F;
            20'd4400: data = 8'h7F;
            20'd4401: data = 8'h7F;
            20'd4402: data = 8'h80;
            20'd4403: data = 8'h80;
            20'd4404: data = 8'h80;
            20'd4405: data = 8'h80;
            20'd4406: data = 8'h80;
            20'd4407: data = 8'h7F;
            20'd4408: data = 8'h80;
            20'd4409: data = 8'h7F;
            20'd4410: data = 8'h7F;
            20'd4411: data = 8'h7F;
            20'd4412: data = 8'h80;
            20'd4413: data = 8'h80;
            20'd4414: data = 8'h80;
            20'd4415: data = 8'h7F;
            20'd4416: data = 8'h80;
            20'd4417: data = 8'h80;
            20'd4418: data = 8'h80;
            20'd4419: data = 8'h80;
            20'd4420: data = 8'h7F;
            20'd4421: data = 8'h80;
            20'd4422: data = 8'h80;
            20'd4423: data = 8'h7F;
            20'd4424: data = 8'h7F;
            20'd4425: data = 8'h80;
            20'd4426: data = 8'h80;
            20'd4427: data = 8'h80;
            20'd4428: data = 8'h7F;
            20'd4429: data = 8'h80;
            20'd4430: data = 8'h80;
            20'd4431: data = 8'h7F;
            20'd4432: data = 8'h7F;
            20'd4433: data = 8'h80;
            20'd4434: data = 8'h80;
            20'd4435: data = 8'h7F;
            20'd4436: data = 8'h80;
            20'd4437: data = 8'h80;
            20'd4438: data = 8'h80;
            20'd4439: data = 8'h80;
            20'd4440: data = 8'h7F;
            20'd4441: data = 8'h7F;
            20'd4442: data = 8'h7F;
            20'd4443: data = 8'h80;
            20'd4444: data = 8'h7F;
            20'd4445: data = 8'h80;
            20'd4446: data = 8'h80;
            20'd4447: data = 8'h80;
            20'd4448: data = 8'h80;
            20'd4449: data = 8'h7F;
            20'd4450: data = 8'h7F;
            20'd4451: data = 8'h80;
            20'd4452: data = 8'h7F;
            20'd4453: data = 8'h80;
            20'd4454: data = 8'h80;
            20'd4455: data = 8'h80;
            20'd4456: data = 8'h7F;
            20'd4457: data = 8'h80;
            20'd4458: data = 8'h80;
            20'd4459: data = 8'h80;
            20'd4460: data = 8'h80;
            20'd4461: data = 8'h7F;
            20'd4462: data = 8'h80;
            20'd4463: data = 8'h80;
            20'd4464: data = 8'h80;
            20'd4465: data = 8'h7F;
            20'd4466: data = 8'h80;
            20'd4467: data = 8'h80;
            20'd4468: data = 8'h80;
            20'd4469: data = 8'h80;
            20'd4470: data = 8'h80;
            20'd4471: data = 8'h7F;
            20'd4472: data = 8'h80;
            20'd4473: data = 8'h80;
            20'd4474: data = 8'h7F;
            20'd4475: data = 8'h7F;
            20'd4476: data = 8'h80;
            20'd4477: data = 8'h80;
            20'd4478: data = 8'h80;
            20'd4479: data = 8'h80;
            20'd4480: data = 8'h80;
            20'd4481: data = 8'h80;
            20'd4482: data = 8'h7F;
            20'd4483: data = 8'h7F;
            20'd4484: data = 8'h80;
            20'd4485: data = 8'h7F;
            20'd4486: data = 8'h80;
            20'd4487: data = 8'h80;
            20'd4488: data = 8'h80;
            20'd4489: data = 8'h7F;
            20'd4490: data = 8'h80;
            20'd4491: data = 8'h7F;
            20'd4492: data = 8'h7F;
            20'd4493: data = 8'h80;
            20'd4494: data = 8'h7F;
            20'd4495: data = 8'h80;
            20'd4496: data = 8'h80;
            20'd4497: data = 8'h7F;
            20'd4498: data = 8'h80;
            20'd4499: data = 8'h80;
            20'd4500: data = 8'h7F;
            20'd4501: data = 8'h80;
            20'd4502: data = 8'h7F;
            20'd4503: data = 8'h7F;
            20'd4504: data = 8'h7F;
            20'd4505: data = 8'h80;
            20'd4506: data = 8'h80;
            20'd4507: data = 8'h80;
            20'd4508: data = 8'h7F;
            20'd4509: data = 8'h80;
            20'd4510: data = 8'h80;
            20'd4511: data = 8'h80;
            20'd4512: data = 8'h80;
            20'd4513: data = 8'h80;
            20'd4514: data = 8'h7F;
            20'd4515: data = 8'h80;
            20'd4516: data = 8'h80;
            20'd4517: data = 8'h80;
            20'd4518: data = 8'h80;
            20'd4519: data = 8'h7F;
            20'd4520: data = 8'h80;
            20'd4521: data = 8'h80;
            20'd4522: data = 8'h80;
            20'd4523: data = 8'h80;
            20'd4524: data = 8'h80;
            20'd4525: data = 8'h80;
            20'd4526: data = 8'h7F;
            20'd4527: data = 8'h80;
            20'd4528: data = 8'h7F;
            20'd4529: data = 8'h80;
            20'd4530: data = 8'h7F;
            20'd4531: data = 8'h80;
            20'd4532: data = 8'h80;
            20'd4533: data = 8'h7F;
            20'd4534: data = 8'h7F;
            20'd4535: data = 8'h80;
            20'd4536: data = 8'h80;
            20'd4537: data = 8'h7F;
            20'd4538: data = 8'h7F;
            20'd4539: data = 8'h80;
            20'd4540: data = 8'h7F;
            20'd4541: data = 8'h7F;
            20'd4542: data = 8'h7F;
            20'd4543: data = 8'h80;
            20'd4544: data = 8'h7F;
            20'd4545: data = 8'h80;
            20'd4546: data = 8'h80;
            20'd4547: data = 8'h7F;
            20'd4548: data = 8'h80;
            20'd4549: data = 8'h80;
            20'd4550: data = 8'h80;
            20'd4551: data = 8'h7F;
            20'd4552: data = 8'h80;
            20'd4553: data = 8'h80;
            20'd4554: data = 8'h80;
            20'd4555: data = 8'h80;
            20'd4556: data = 8'h80;
            20'd4557: data = 8'h80;
            20'd4558: data = 8'h80;
            20'd4559: data = 8'h80;
            20'd4560: data = 8'h80;
            20'd4561: data = 8'h80;
            20'd4562: data = 8'h80;
            20'd4563: data = 8'h80;
            20'd4564: data = 8'h80;
            20'd4565: data = 8'h7F;
            20'd4566: data = 8'h80;
            20'd4567: data = 8'h80;
            20'd4568: data = 8'h80;
            20'd4569: data = 8'h80;
            20'd4570: data = 8'h7F;
            20'd4571: data = 8'h80;
            20'd4572: data = 8'h80;
            20'd4573: data = 8'h7F;
            20'd4574: data = 8'h80;
            20'd4575: data = 8'h80;
            20'd4576: data = 8'h7F;
            20'd4577: data = 8'h7F;
            20'd4578: data = 8'h7F;
            20'd4579: data = 8'h80;
            20'd4580: data = 8'h7F;
            20'd4581: data = 8'h80;
            20'd4582: data = 8'h80;
            20'd4583: data = 8'h7F;
            20'd4584: data = 8'h7F;
            20'd4585: data = 8'h80;
            20'd4586: data = 8'h80;
            20'd4587: data = 8'h7F;
            20'd4588: data = 8'h80;
            20'd4589: data = 8'h7F;
            20'd4590: data = 8'h80;
            20'd4591: data = 8'h80;
            20'd4592: data = 8'h80;
            20'd4593: data = 8'h80;
            20'd4594: data = 8'h80;
            20'd4595: data = 8'h80;
            20'd4596: data = 8'h80;
            20'd4597: data = 8'h7F;
            20'd4598: data = 8'h80;
            20'd4599: data = 8'h80;
            20'd4600: data = 8'h7F;
            20'd4601: data = 8'h80;
            20'd4602: data = 8'h80;
            20'd4603: data = 8'h80;
            20'd4604: data = 8'h80;
            20'd4605: data = 8'h80;
            20'd4606: data = 8'h80;
            20'd4607: data = 8'h80;
            20'd4608: data = 8'h80;
            20'd4609: data = 8'h7F;
            20'd4610: data = 8'h80;
            20'd4611: data = 8'h80;
            20'd4612: data = 8'h80;
            20'd4613: data = 8'h80;
            20'd4614: data = 8'h7F;
            20'd4615: data = 8'h7F;
            20'd4616: data = 8'h7F;
            20'd4617: data = 8'h7F;
            20'd4618: data = 8'h80;
            20'd4619: data = 8'h80;
            20'd4620: data = 8'h80;
            20'd4621: data = 8'h80;
            20'd4622: data = 8'h80;
            20'd4623: data = 8'h80;
            20'd4624: data = 8'h80;
            20'd4625: data = 8'h7F;
            20'd4626: data = 8'h80;
            20'd4627: data = 8'h80;
            20'd4628: data = 8'h80;
            20'd4629: data = 8'h80;
            20'd4630: data = 8'h7F;
            20'd4631: data = 8'h80;
            20'd4632: data = 8'h80;
            20'd4633: data = 8'h80;
            20'd4634: data = 8'h80;
            20'd4635: data = 8'h7F;
            20'd4636: data = 8'h7F;
            20'd4637: data = 8'h7F;
            20'd4638: data = 8'h80;
            20'd4639: data = 8'h80;
            20'd4640: data = 8'h80;
            20'd4641: data = 8'h80;
            20'd4642: data = 8'h80;
            20'd4643: data = 8'h7F;
            20'd4644: data = 8'h7F;
            20'd4645: data = 8'h80;
            20'd4646: data = 8'h80;
            20'd4647: data = 8'h80;
            20'd4648: data = 8'h80;
            20'd4649: data = 8'h7F;
            20'd4650: data = 8'h80;
            20'd4651: data = 8'h80;
            20'd4652: data = 8'h7F;
            20'd4653: data = 8'h80;
            20'd4654: data = 8'h80;
            20'd4655: data = 8'h80;
            20'd4656: data = 8'h80;
            20'd4657: data = 8'h7F;
            20'd4658: data = 8'h7F;
            20'd4659: data = 8'h80;
            20'd4660: data = 8'h80;
            20'd4661: data = 8'h80;
            20'd4662: data = 8'h80;
            20'd4663: data = 8'h7F;
            20'd4664: data = 8'h80;
            20'd4665: data = 8'h7F;
            20'd4666: data = 8'h80;
            20'd4667: data = 8'h80;
            20'd4668: data = 8'h80;
            20'd4669: data = 8'h80;
            20'd4670: data = 8'h7F;
            20'd4671: data = 8'h80;
            20'd4672: data = 8'h80;
            20'd4673: data = 8'h80;
            20'd4674: data = 8'h7F;
            20'd4675: data = 8'h80;
            20'd4676: data = 8'h80;
            20'd4677: data = 8'h80;
            20'd4678: data = 8'h7F;
            20'd4679: data = 8'h80;
            20'd4680: data = 8'h7F;
            20'd4681: data = 8'h7F;
            20'd4682: data = 8'h80;
            20'd4683: data = 8'h7F;
            20'd4684: data = 8'h80;
            20'd4685: data = 8'h80;
            20'd4686: data = 8'h7F;
            20'd4687: data = 8'h7F;
            20'd4688: data = 8'h80;
            20'd4689: data = 8'h80;
            20'd4690: data = 8'h7F;
            20'd4691: data = 8'h80;
            20'd4692: data = 8'h7F;
            20'd4693: data = 8'h7F;
            20'd4694: data = 8'h80;
            20'd4695: data = 8'h80;
            20'd4696: data = 8'h80;
            20'd4697: data = 8'h80;
            20'd4698: data = 8'h80;
            20'd4699: data = 8'h80;
            20'd4700: data = 8'h80;
            20'd4701: data = 8'h80;
            20'd4702: data = 8'h80;
            20'd4703: data = 8'h7F;
            20'd4704: data = 8'h7F;
            20'd4705: data = 8'h80;
            20'd4706: data = 8'h7F;
            20'd4707: data = 8'h80;
            20'd4708: data = 8'h7F;
            20'd4709: data = 8'h80;
            20'd4710: data = 8'h80;
            20'd4711: data = 8'h80;
            20'd4712: data = 8'h7F;
            20'd4713: data = 8'h80;
            20'd4714: data = 8'h80;
            20'd4715: data = 8'h7F;
            20'd4716: data = 8'h80;
            20'd4717: data = 8'h80;
            20'd4718: data = 8'h7F;
            20'd4719: data = 8'h7F;
            20'd4720: data = 8'h80;
            20'd4721: data = 8'h80;
            20'd4722: data = 8'h80;
            20'd4723: data = 8'h7F;
            20'd4724: data = 8'h80;
            20'd4725: data = 8'h80;
            20'd4726: data = 8'h80;
            20'd4727: data = 8'h80;
            20'd4728: data = 8'h80;
            20'd4729: data = 8'h7F;
            20'd4730: data = 8'h80;
            20'd4731: data = 8'h7F;
            20'd4732: data = 8'h80;
            20'd4733: data = 8'h80;
            20'd4734: data = 8'h7F;
            20'd4735: data = 8'h80;
            20'd4736: data = 8'h80;
            20'd4737: data = 8'h80;
            20'd4738: data = 8'h80;
            20'd4739: data = 8'h7F;
            20'd4740: data = 8'h7F;
            20'd4741: data = 8'h80;
            20'd4742: data = 8'h80;
            20'd4743: data = 8'h80;
            20'd4744: data = 8'h80;
            20'd4745: data = 8'h80;
            20'd4746: data = 8'h80;
            20'd4747: data = 8'h7F;
            20'd4748: data = 8'h80;
            20'd4749: data = 8'h80;
            20'd4750: data = 8'h7F;
            20'd4751: data = 8'h80;
            20'd4752: data = 8'h80;
            20'd4753: data = 8'h80;
            20'd4754: data = 8'h7F;
            20'd4755: data = 8'h80;
            20'd4756: data = 8'h80;
            20'd4757: data = 8'h7F;
            20'd4758: data = 8'h7F;
            20'd4759: data = 8'h80;
            20'd4760: data = 8'h80;
            20'd4761: data = 8'h80;
            20'd4762: data = 8'h80;
            20'd4763: data = 8'h80;
            20'd4764: data = 8'h80;
            20'd4765: data = 8'h7F;
            20'd4766: data = 8'h80;
            20'd4767: data = 8'h80;
            20'd4768: data = 8'h80;
            20'd4769: data = 8'h80;
            20'd4770: data = 8'h80;
            20'd4771: data = 8'h80;
            20'd4772: data = 8'h80;
            20'd4773: data = 8'h80;
            20'd4774: data = 8'h7F;
            20'd4775: data = 8'h80;
            20'd4776: data = 8'h80;
            20'd4777: data = 8'h7F;
            20'd4778: data = 8'h80;
            20'd4779: data = 8'h80;
            20'd4780: data = 8'h80;
            20'd4781: data = 8'h7F;
            20'd4782: data = 8'h80;
            20'd4783: data = 8'h80;
            20'd4784: data = 8'h80;
            20'd4785: data = 8'h80;
            20'd4786: data = 8'h7F;
            20'd4787: data = 8'h7F;
            20'd4788: data = 8'h80;
            20'd4789: data = 8'h80;
            20'd4790: data = 8'h80;
            20'd4791: data = 8'h80;
            20'd4792: data = 8'h80;
            20'd4793: data = 8'h80;
            20'd4794: data = 8'h7F;
            20'd4795: data = 8'h7F;
            20'd4796: data = 8'h80;
            20'd4797: data = 8'h80;
            20'd4798: data = 8'h80;
            20'd4799: data = 8'h80;
            20'd4800: data = 8'h80;
            20'd4801: data = 8'h80;
            20'd4802: data = 8'h80;
            20'd4803: data = 8'h7F;
            20'd4804: data = 8'h80;
            20'd4805: data = 8'h7F;
            20'd4806: data = 8'h7F;
            20'd4807: data = 8'h80;
            20'd4808: data = 8'h80;
            20'd4809: data = 8'h80;
            20'd4810: data = 8'h80;
            20'd4811: data = 8'h7F;
            20'd4812: data = 8'h7F;
            20'd4813: data = 8'h80;
            20'd4814: data = 8'h80;
            20'd4815: data = 8'h80;
            20'd4816: data = 8'h80;
            20'd4817: data = 8'h80;
            20'd4818: data = 8'h80;
            20'd4819: data = 8'h80;
            20'd4820: data = 8'h7F;
            20'd4821: data = 8'h80;
            20'd4822: data = 8'h7F;
            20'd4823: data = 8'h80;
            20'd4824: data = 8'h80;
            20'd4825: data = 8'h80;
            20'd4826: data = 8'h7F;
            20'd4827: data = 8'h7F;
            20'd4828: data = 8'h80;
            20'd4829: data = 8'h80;
            20'd4830: data = 8'h7F;
            20'd4831: data = 8'h80;
            20'd4832: data = 8'h7F;
            20'd4833: data = 8'h80;
            20'd4834: data = 8'h80;
            20'd4835: data = 8'h80;
            20'd4836: data = 8'h7F;
            20'd4837: data = 8'h80;
            20'd4838: data = 8'h7F;
            20'd4839: data = 8'h7F;
            20'd4840: data = 8'h7F;
            20'd4841: data = 8'h80;
            20'd4842: data = 8'h7F;
            20'd4843: data = 8'h80;
            20'd4844: data = 8'h80;
            20'd4845: data = 8'h80;
            20'd4846: data = 8'h80;
            20'd4847: data = 8'h80;
            20'd4848: data = 8'h80;
            20'd4849: data = 8'h7F;
            20'd4850: data = 8'h80;
            20'd4851: data = 8'h7F;
            20'd4852: data = 8'h80;
            20'd4853: data = 8'h7F;
            20'd4854: data = 8'h80;
            20'd4855: data = 8'h80;
            20'd4856: data = 8'h80;
            20'd4857: data = 8'h7F;
            20'd4858: data = 8'h7F;
            20'd4859: data = 8'h80;
            20'd4860: data = 8'h7F;
            20'd4861: data = 8'h7F;
            20'd4862: data = 8'h80;
            20'd4863: data = 8'h80;
            20'd4864: data = 8'h80;
            20'd4865: data = 8'h80;
            20'd4866: data = 8'h80;
            20'd4867: data = 8'h80;
            20'd4868: data = 8'h80;
            20'd4869: data = 8'h80;
            20'd4870: data = 8'h80;
            20'd4871: data = 8'h80;
            20'd4872: data = 8'h80;
            20'd4873: data = 8'h80;
            20'd4874: data = 8'h7F;
            20'd4875: data = 8'h7F;
            20'd4876: data = 8'h7F;
            20'd4877: data = 8'h80;
            20'd4878: data = 8'h80;
            20'd4879: data = 8'h80;
            20'd4880: data = 8'h7F;
            20'd4881: data = 8'h7F;
            20'd4882: data = 8'h80;
            20'd4883: data = 8'h80;
            20'd4884: data = 8'h7F;
            20'd4885: data = 8'h7F;
            20'd4886: data = 8'h80;
            20'd4887: data = 8'h80;
            20'd4888: data = 8'h7F;
            20'd4889: data = 8'h7F;
            20'd4890: data = 8'h80;
            20'd4891: data = 8'h80;
            20'd4892: data = 8'h80;
            20'd4893: data = 8'h80;
            20'd4894: data = 8'h7F;
            20'd4895: data = 8'h7F;
            20'd4896: data = 8'h80;
            20'd4897: data = 8'h80;
            20'd4898: data = 8'h80;
            20'd4899: data = 8'h80;
            20'd4900: data = 8'h7F;
            20'd4901: data = 8'h80;
            20'd4902: data = 8'h80;
            20'd4903: data = 8'h7F;
            20'd4904: data = 8'h80;
            20'd4905: data = 8'h80;
            20'd4906: data = 8'h80;
            20'd4907: data = 8'h7F;
            20'd4908: data = 8'h7F;
            20'd4909: data = 8'h7F;
            20'd4910: data = 8'h7F;
            20'd4911: data = 8'h80;
            20'd4912: data = 8'h80;
            20'd4913: data = 8'h80;
            20'd4914: data = 8'h80;
            20'd4915: data = 8'h80;
            20'd4916: data = 8'h7F;
            20'd4917: data = 8'h80;
            20'd4918: data = 8'h80;
            20'd4919: data = 8'h80;
            20'd4920: data = 8'h7F;
            20'd4921: data = 8'h80;
            20'd4922: data = 8'h80;
            20'd4923: data = 8'h80;
            20'd4924: data = 8'h80;
            20'd4925: data = 8'h80;
            20'd4926: data = 8'h80;
            20'd4927: data = 8'h80;
            20'd4928: data = 8'h7F;
            20'd4929: data = 8'h80;
            20'd4930: data = 8'h80;
            20'd4931: data = 8'h80;
            20'd4932: data = 8'h7F;
            20'd4933: data = 8'h80;
            20'd4934: data = 8'h7F;
            20'd4935: data = 8'h7F;
            20'd4936: data = 8'h80;
            20'd4937: data = 8'h80;
            20'd4938: data = 8'h80;
            20'd4939: data = 8'h80;
            20'd4940: data = 8'h7F;
            20'd4941: data = 8'h80;
            20'd4942: data = 8'h80;
            20'd4943: data = 8'h80;
            20'd4944: data = 8'h80;
            20'd4945: data = 8'h7F;
            20'd4946: data = 8'h7F;
            20'd4947: data = 8'h80;
            20'd4948: data = 8'h7F;
            20'd4949: data = 8'h80;
            20'd4950: data = 8'h7F;
            20'd4951: data = 8'h7F;
            20'd4952: data = 8'h7F;
            20'd4953: data = 8'h80;
            20'd4954: data = 8'h7F;
            20'd4955: data = 8'h80;
            20'd4956: data = 8'h80;
            20'd4957: data = 8'h80;
            20'd4958: data = 8'h80;
            20'd4959: data = 8'h7F;
            20'd4960: data = 8'h7F;
            20'd4961: data = 8'h80;
            20'd4962: data = 8'h80;
            20'd4963: data = 8'h7F;
            20'd4964: data = 8'h80;
            20'd4965: data = 8'h80;
            20'd4966: data = 8'h80;
            20'd4967: data = 8'h80;
            20'd4968: data = 8'h80;
            20'd4969: data = 8'h7F;
            20'd4970: data = 8'h80;
            20'd4971: data = 8'h80;
            20'd4972: data = 8'h7F;
            20'd4973: data = 8'h80;
            20'd4974: data = 8'h80;
            20'd4975: data = 8'h80;
            20'd4976: data = 8'h80;
            20'd4977: data = 8'h80;
            20'd4978: data = 8'h80;
            20'd4979: data = 8'h80;
            20'd4980: data = 8'h7F;
            20'd4981: data = 8'h7F;
            20'd4982: data = 8'h80;
            20'd4983: data = 8'h80;
            20'd4984: data = 8'h80;
            20'd4985: data = 8'h7F;
            20'd4986: data = 8'h80;
            20'd4987: data = 8'h80;
            20'd4988: data = 8'h80;
            20'd4989: data = 8'h80;
            20'd4990: data = 8'h80;
            20'd4991: data = 8'h7F;
            20'd4992: data = 8'h80;
            20'd4993: data = 8'h80;
            20'd4994: data = 8'h80;
            20'd4995: data = 8'h7F;
            20'd4996: data = 8'h80;
            20'd4997: data = 8'h80;
            20'd4998: data = 8'h7F;
            20'd4999: data = 8'h80;
            20'd5000: data = 8'h80;
            20'd5001: data = 8'h7F;
            20'd5002: data = 8'h80;
            20'd5003: data = 8'h80;
            20'd5004: data = 8'h7F;
            20'd5005: data = 8'h7F;
            20'd5006: data = 8'h7F;
            20'd5007: data = 8'h80;
            20'd5008: data = 8'h80;
            20'd5009: data = 8'h7F;
            20'd5010: data = 8'h80;
            20'd5011: data = 8'h80;
            20'd5012: data = 8'h80;
            20'd5013: data = 8'h7F;
            20'd5014: data = 8'h7F;
            20'd5015: data = 8'h80;
            20'd5016: data = 8'h80;
            20'd5017: data = 8'h7F;
            20'd5018: data = 8'h80;
            20'd5019: data = 8'h80;
            20'd5020: data = 8'h80;
            20'd5021: data = 8'h7F;
            20'd5022: data = 8'h7F;
            20'd5023: data = 8'h80;
            20'd5024: data = 8'h80;
            20'd5025: data = 8'h7F;
            20'd5026: data = 8'h80;
            20'd5027: data = 8'h80;
            20'd5028: data = 8'h80;
            20'd5029: data = 8'h7F;
            20'd5030: data = 8'h7F;
            20'd5031: data = 8'h80;
            20'd5032: data = 8'h80;
            20'd5033: data = 8'h80;
            20'd5034: data = 8'h80;
            20'd5035: data = 8'h7F;
            20'd5036: data = 8'h80;
            20'd5037: data = 8'h80;
            20'd5038: data = 8'h80;
            20'd5039: data = 8'h80;
            20'd5040: data = 8'h80;
            20'd5041: data = 8'h80;
            20'd5042: data = 8'h80;
            20'd5043: data = 8'h7F;
            20'd5044: data = 8'h80;
            20'd5045: data = 8'h80;
            20'd5046: data = 8'h80;
            20'd5047: data = 8'h80;
            20'd5048: data = 8'h80;
            20'd5049: data = 8'h80;
            20'd5050: data = 8'h80;
            20'd5051: data = 8'h7F;
            20'd5052: data = 8'h80;
            20'd5053: data = 8'h80;
            20'd5054: data = 8'h80;
            20'd5055: data = 8'h7F;
            20'd5056: data = 8'h7F;
            20'd5057: data = 8'h80;
            20'd5058: data = 8'h80;
            20'd5059: data = 8'h7F;
            20'd5060: data = 8'h7F;
            20'd5061: data = 8'h80;
            20'd5062: data = 8'h80;
            20'd5063: data = 8'h80;
            20'd5064: data = 8'h80;
            20'd5065: data = 8'h7F;
            20'd5066: data = 8'h80;
            20'd5067: data = 8'h80;
            20'd5068: data = 8'h80;
            20'd5069: data = 8'h80;
            20'd5070: data = 8'h80;
            20'd5071: data = 8'h80;
            20'd5072: data = 8'h80;
            20'd5073: data = 8'h80;
            20'd5074: data = 8'h80;
            20'd5075: data = 8'h80;
            20'd5076: data = 8'h80;
            20'd5077: data = 8'h7F;
            20'd5078: data = 8'h80;
            20'd5079: data = 8'h80;
            20'd5080: data = 8'h80;
            20'd5081: data = 8'h80;
            20'd5082: data = 8'h7F;
            20'd5083: data = 8'h7F;
            20'd5084: data = 8'h80;
            20'd5085: data = 8'h80;
            20'd5086: data = 8'h7F;
            20'd5087: data = 8'h80;
            20'd5088: data = 8'h7F;
            20'd5089: data = 8'h80;
            20'd5090: data = 8'h7F;
            20'd5091: data = 8'h80;
            20'd5092: data = 8'h80;
            20'd5093: data = 8'h7F;
            20'd5094: data = 8'h80;
            20'd5095: data = 8'h7F;
            20'd5096: data = 8'h80;
            20'd5097: data = 8'h80;
            20'd5098: data = 8'h7F;
            20'd5099: data = 8'h7F;
            20'd5100: data = 8'h7F;
            20'd5101: data = 8'h80;
            20'd5102: data = 8'h7F;
            20'd5103: data = 8'h80;
            20'd5104: data = 8'h80;
            20'd5105: data = 8'h7F;
            20'd5106: data = 8'h7F;
            20'd5107: data = 8'h80;
            20'd5108: data = 8'h80;
            20'd5109: data = 8'h80;
            20'd5110: data = 8'h80;
            20'd5111: data = 8'h80;
            20'd5112: data = 8'h80;
            20'd5113: data = 8'h80;
            20'd5114: data = 8'h80;
            20'd5115: data = 8'h7F;
            20'd5116: data = 8'h80;
            20'd5117: data = 8'h80;
            20'd5118: data = 8'h80;
            20'd5119: data = 8'h7F;
            20'd5120: data = 8'h80;
            20'd5121: data = 8'h80;
            20'd5122: data = 8'h7F;
            20'd5123: data = 8'h7F;
            20'd5124: data = 8'h80;
            20'd5125: data = 8'h80;
            20'd5126: data = 8'h7F;
            20'd5127: data = 8'h80;
            20'd5128: data = 8'h80;
            20'd5129: data = 8'h80;
            20'd5130: data = 8'h7F;
            20'd5131: data = 8'h80;
            20'd5132: data = 8'h80;
            20'd5133: data = 8'h7F;
            20'd5134: data = 8'h7F;
            20'd5135: data = 8'h80;
            20'd5136: data = 8'h80;
            20'd5137: data = 8'h80;
            20'd5138: data = 8'h80;
            20'd5139: data = 8'h80;
            20'd5140: data = 8'h7F;
            20'd5141: data = 8'h80;
            20'd5142: data = 8'h80;
            20'd5143: data = 8'h80;
            20'd5144: data = 8'h7F;
            20'd5145: data = 8'h80;
            20'd5146: data = 8'h80;
            20'd5147: data = 8'h80;
            20'd5148: data = 8'h80;
            20'd5149: data = 8'h80;
            20'd5150: data = 8'h80;
            20'd5151: data = 8'h80;
            20'd5152: data = 8'h80;
            20'd5153: data = 8'h80;
            20'd5154: data = 8'h80;
            20'd5155: data = 8'h80;
            20'd5156: data = 8'h80;
            20'd5157: data = 8'h7F;
            20'd5158: data = 8'h7F;
            20'd5159: data = 8'h80;
            20'd5160: data = 8'h80;
            20'd5161: data = 8'h80;
            20'd5162: data = 8'h80;
            20'd5163: data = 8'h80;
            20'd5164: data = 8'h7F;
            20'd5165: data = 8'h80;
            20'd5166: data = 8'h80;
            20'd5167: data = 8'h80;
            20'd5168: data = 8'h7F;
            20'd5169: data = 8'h80;
            20'd5170: data = 8'h80;
            20'd5171: data = 8'h80;
            20'd5172: data = 8'h80;
            20'd5173: data = 8'h80;
            20'd5174: data = 8'h80;
            20'd5175: data = 8'h7F;
            20'd5176: data = 8'h80;
            20'd5177: data = 8'h7F;
            20'd5178: data = 8'h80;
            20'd5179: data = 8'h80;
            20'd5180: data = 8'h80;
            20'd5181: data = 8'h7F;
            20'd5182: data = 8'h80;
            20'd5183: data = 8'h80;
            20'd5184: data = 8'h80;
            20'd5185: data = 8'h7F;
            20'd5186: data = 8'h80;
            20'd5187: data = 8'h80;
            20'd5188: data = 8'h80;
            20'd5189: data = 8'h80;
            20'd5190: data = 8'h80;
            20'd5191: data = 8'h7F;
            20'd5192: data = 8'h80;
            20'd5193: data = 8'h7F;
            20'd5194: data = 8'h80;
            20'd5195: data = 8'h80;
            20'd5196: data = 8'h7F;
            20'd5197: data = 8'h80;
            20'd5198: data = 8'h80;
            20'd5199: data = 8'h7F;
            20'd5200: data = 8'h80;
            20'd5201: data = 8'h7F;
            20'd5202: data = 8'h7F;
            20'd5203: data = 8'h80;
            20'd5204: data = 8'h7F;
            20'd5205: data = 8'h7F;
            20'd5206: data = 8'h80;
            20'd5207: data = 8'h80;
            20'd5208: data = 8'h7F;
            20'd5209: data = 8'h7F;
            20'd5210: data = 8'h80;
            20'd5211: data = 8'h7F;
            20'd5212: data = 8'h80;
            20'd5213: data = 8'h80;
            20'd5214: data = 8'h7F;
            20'd5215: data = 8'h7F;
            20'd5216: data = 8'h80;
            20'd5217: data = 8'h7F;
            20'd5218: data = 8'h80;
            20'd5219: data = 8'h7F;
            20'd5220: data = 8'h7F;
            20'd5221: data = 8'h80;
            20'd5222: data = 8'h80;
            20'd5223: data = 8'h7F;
            20'd5224: data = 8'h7F;
            20'd5225: data = 8'h7F;
            20'd5226: data = 8'h80;
            20'd5227: data = 8'h80;
            20'd5228: data = 8'h7F;
            20'd5229: data = 8'h80;
            20'd5230: data = 8'h80;
            20'd5231: data = 8'h7F;
            20'd5232: data = 8'h7F;
            20'd5233: data = 8'h80;
            20'd5234: data = 8'h80;
            20'd5235: data = 8'h80;
            20'd5236: data = 8'h7F;
            20'd5237: data = 8'h7F;
            20'd5238: data = 8'h80;
            20'd5239: data = 8'h80;
            20'd5240: data = 8'h7F;
            20'd5241: data = 8'h80;
            20'd5242: data = 8'h7F;
            20'd5243: data = 8'h80;
            20'd5244: data = 8'h80;
            20'd5245: data = 8'h80;
            20'd5246: data = 8'h80;
            20'd5247: data = 8'h7F;
            20'd5248: data = 8'h80;
            20'd5249: data = 8'h7F;
            20'd5250: data = 8'h7F;
            20'd5251: data = 8'h80;
            20'd5252: data = 8'h80;
            20'd5253: data = 8'h7F;
            20'd5254: data = 8'h7F;
            20'd5255: data = 8'h80;
            20'd5256: data = 8'h80;
            20'd5257: data = 8'h80;
            20'd5258: data = 8'h7F;
            20'd5259: data = 8'h80;
            20'd5260: data = 8'h7F;
            20'd5261: data = 8'h7F;
            20'd5262: data = 8'h80;
            20'd5263: data = 8'h80;
            20'd5264: data = 8'h7F;
            20'd5265: data = 8'h7F;
            20'd5266: data = 8'h80;
            20'd5267: data = 8'h80;
            20'd5268: data = 8'h7F;
            20'd5269: data = 8'h7F;
            20'd5270: data = 8'h80;
            20'd5271: data = 8'h7F;
            20'd5272: data = 8'h7F;
            20'd5273: data = 8'h80;
            20'd5274: data = 8'h80;
            20'd5275: data = 8'h80;
            20'd5276: data = 8'h80;
            20'd5277: data = 8'h7F;
            20'd5278: data = 8'h7F;
            20'd5279: data = 8'h80;
            20'd5280: data = 8'h7F;
            20'd5281: data = 8'h7F;
            20'd5282: data = 8'h80;
            20'd5283: data = 8'h80;
            20'd5284: data = 8'h7F;
            20'd5285: data = 8'h7F;
            20'd5286: data = 8'h80;
            20'd5287: data = 8'h7F;
            20'd5288: data = 8'h80;
            20'd5289: data = 8'h80;
            20'd5290: data = 8'h80;
            20'd5291: data = 8'h80;
            20'd5292: data = 8'h7F;
            20'd5293: data = 8'h80;
            20'd5294: data = 8'h80;
            20'd5295: data = 8'h80;
            20'd5296: data = 8'h80;
            20'd5297: data = 8'h80;
            20'd5298: data = 8'h7F;
            20'd5299: data = 8'h80;
            20'd5300: data = 8'h80;
            20'd5301: data = 8'h80;
            20'd5302: data = 8'h80;
            20'd5303: data = 8'h80;
            20'd5304: data = 8'h80;
            20'd5305: data = 8'h80;
            20'd5306: data = 8'h7F;
            20'd5307: data = 8'h7F;
            20'd5308: data = 8'h80;
            20'd5309: data = 8'h80;
            20'd5310: data = 8'h80;
            20'd5311: data = 8'h7F;
            20'd5312: data = 8'h7F;
            20'd5313: data = 8'h80;
            20'd5314: data = 8'h80;
            20'd5315: data = 8'h80;
            20'd5316: data = 8'h80;
            20'd5317: data = 8'h7F;
            20'd5318: data = 8'h7F;
            20'd5319: data = 8'h80;
            20'd5320: data = 8'h80;
            20'd5321: data = 8'h80;
            20'd5322: data = 8'h7F;
            20'd5323: data = 8'h80;
            20'd5324: data = 8'h80;
            20'd5325: data = 8'h7F;
            20'd5326: data = 8'h80;
            20'd5327: data = 8'h80;
            20'd5328: data = 8'h80;
            20'd5329: data = 8'h80;
            20'd5330: data = 8'h7F;
            20'd5331: data = 8'h80;
            20'd5332: data = 8'h80;
            20'd5333: data = 8'h7F;
            20'd5334: data = 8'h7F;
            20'd5335: data = 8'h80;
            20'd5336: data = 8'h7F;
            20'd5337: data = 8'h7F;
            20'd5338: data = 8'h7F;
            20'd5339: data = 8'h80;
            20'd5340: data = 8'h80;
            20'd5341: data = 8'h7F;
            20'd5342: data = 8'h7F;
            20'd5343: data = 8'h80;
            20'd5344: data = 8'h7F;
            20'd5345: data = 8'h7F;
            20'd5346: data = 8'h80;
            20'd5347: data = 8'h7F;
            20'd5348: data = 8'h80;
            20'd5349: data = 8'h80;
            20'd5350: data = 8'h80;
            20'd5351: data = 8'h7F;
            20'd5352: data = 8'h7F;
            20'd5353: data = 8'h7F;
            20'd5354: data = 8'h80;
            20'd5355: data = 8'h80;
            20'd5356: data = 8'h80;
            20'd5357: data = 8'h80;
            20'd5358: data = 8'h80;
            20'd5359: data = 8'h80;
            20'd5360: data = 8'h80;
            20'd5361: data = 8'h7F;
            20'd5362: data = 8'h80;
            20'd5363: data = 8'h7F;
            20'd5364: data = 8'h7F;
            20'd5365: data = 8'h80;
            20'd5366: data = 8'h80;
            20'd5367: data = 8'h80;
            20'd5368: data = 8'h80;
            20'd5369: data = 8'h80;
            20'd5370: data = 8'h7F;
            20'd5371: data = 8'h80;
            20'd5372: data = 8'h80;
            20'd5373: data = 8'h80;
            20'd5374: data = 8'h7F;
            20'd5375: data = 8'h80;
            20'd5376: data = 8'h80;
            20'd5377: data = 8'h80;
            20'd5378: data = 8'h80;
            20'd5379: data = 8'h80;
            20'd5380: data = 8'h80;
            20'd5381: data = 8'h80;
            20'd5382: data = 8'h7F;
            20'd5383: data = 8'h80;
            20'd5384: data = 8'h80;
            20'd5385: data = 8'h7F;
            20'd5386: data = 8'h7F;
            20'd5387: data = 8'h80;
            20'd5388: data = 8'h80;
            20'd5389: data = 8'h7F;
            20'd5390: data = 8'h7F;
            20'd5391: data = 8'h80;
            20'd5392: data = 8'h80;
            20'd5393: data = 8'h80;
            20'd5394: data = 8'h80;
            20'd5395: data = 8'h7F;
            20'd5396: data = 8'h80;
            20'd5397: data = 8'h80;
            20'd5398: data = 8'h7F;
            20'd5399: data = 8'h80;
            20'd5400: data = 8'h80;
            20'd5401: data = 8'h80;
            20'd5402: data = 8'h80;
            20'd5403: data = 8'h80;
            20'd5404: data = 8'h7F;
            20'd5405: data = 8'h7F;
            20'd5406: data = 8'h80;
            20'd5407: data = 8'h80;
            20'd5408: data = 8'h80;
            20'd5409: data = 8'h80;
            20'd5410: data = 8'h80;
            20'd5411: data = 8'h7F;
            20'd5412: data = 8'h80;
            20'd5413: data = 8'h80;
            20'd5414: data = 8'h80;
            20'd5415: data = 8'h80;
            20'd5416: data = 8'h80;
            20'd5417: data = 8'h7F;
            20'd5418: data = 8'h7F;
            20'd5419: data = 8'h7F;
            20'd5420: data = 8'h80;
            20'd5421: data = 8'h80;
            20'd5422: data = 8'h80;
            20'd5423: data = 8'h7F;
            20'd5424: data = 8'h80;
            20'd5425: data = 8'h80;
            20'd5426: data = 8'h80;
            20'd5427: data = 8'h80;
            20'd5428: data = 8'h80;
            20'd5429: data = 8'h80;
            20'd5430: data = 8'h7F;
            20'd5431: data = 8'h80;
            20'd5432: data = 8'h7F;
            20'd5433: data = 8'h7F;
            20'd5434: data = 8'h80;
            20'd5435: data = 8'h7F;
            20'd5436: data = 8'h80;
            20'd5437: data = 8'h80;
            20'd5438: data = 8'h7F;
            20'd5439: data = 8'h80;
            20'd5440: data = 8'h80;
            20'd5441: data = 8'h7F;
            20'd5442: data = 8'h80;
            20'd5443: data = 8'h80;
            20'd5444: data = 8'h80;
            20'd5445: data = 8'h7F;
            20'd5446: data = 8'h80;
            20'd5447: data = 8'h7F;
            20'd5448: data = 8'h80;
            20'd5449: data = 8'h80;
            20'd5450: data = 8'h80;
            20'd5451: data = 8'h80;
            20'd5452: data = 8'h7F;
            20'd5453: data = 8'h7F;
            20'd5454: data = 8'h7F;
            20'd5455: data = 8'h7F;
            20'd5456: data = 8'h80;
            20'd5457: data = 8'h80;
            20'd5458: data = 8'h80;
            20'd5459: data = 8'h80;
            20'd5460: data = 8'h80;
            20'd5461: data = 8'h80;
            20'd5462: data = 8'h80;
            20'd5463: data = 8'h80;
            20'd5464: data = 8'h7F;
            20'd5465: data = 8'h80;
            20'd5466: data = 8'h7F;
            20'd5467: data = 8'h80;
            20'd5468: data = 8'h7F;
            20'd5469: data = 8'h80;
            20'd5470: data = 8'h7F;
            20'd5471: data = 8'h80;
            20'd5472: data = 8'h80;
            20'd5473: data = 8'h80;
            20'd5474: data = 8'h7F;
            20'd5475: data = 8'h7F;
            20'd5476: data = 8'h80;
            20'd5477: data = 8'h7F;
            20'd5478: data = 8'h80;
            20'd5479: data = 8'h7F;
            20'd5480: data = 8'h80;
            20'd5481: data = 8'h7F;
            20'd5482: data = 8'h7F;
            20'd5483: data = 8'h80;
            20'd5484: data = 8'h7F;
            20'd5485: data = 8'h80;
            20'd5486: data = 8'h80;
            20'd5487: data = 8'h80;
            20'd5488: data = 8'h80;
            20'd5489: data = 8'h7F;
            20'd5490: data = 8'h80;
            20'd5491: data = 8'h80;
            20'd5492: data = 8'h80;
            20'd5493: data = 8'h80;
            20'd5494: data = 8'h7F;
            20'd5495: data = 8'h80;
            20'd5496: data = 8'h80;
            20'd5497: data = 8'h80;
            20'd5498: data = 8'h80;
            20'd5499: data = 8'h80;
            20'd5500: data = 8'h80;
            20'd5501: data = 8'h80;
            20'd5502: data = 8'h80;
            20'd5503: data = 8'h80;
            20'd5504: data = 8'h7F;
            20'd5505: data = 8'h80;
            20'd5506: data = 8'h80;
            20'd5507: data = 8'h80;
            20'd5508: data = 8'h80;
            20'd5509: data = 8'h80;
            20'd5510: data = 8'h80;
            20'd5511: data = 8'h7F;
            20'd5512: data = 8'h7F;
            20'd5513: data = 8'h7F;
            20'd5514: data = 8'h7F;
            20'd5515: data = 8'h80;
            20'd5516: data = 8'h80;
            20'd5517: data = 8'h80;
            20'd5518: data = 8'h7F;
            20'd5519: data = 8'h80;
            20'd5520: data = 8'h80;
            20'd5521: data = 8'h80;
            20'd5522: data = 8'h80;
            20'd5523: data = 8'h80;
            20'd5524: data = 8'h80;
            20'd5525: data = 8'h80;
            20'd5526: data = 8'h80;
            20'd5527: data = 8'h80;
            20'd5528: data = 8'h7F;
            20'd5529: data = 8'h80;
            20'd5530: data = 8'h80;
            20'd5531: data = 8'h80;
            20'd5532: data = 8'h80;
            20'd5533: data = 8'h80;
            20'd5534: data = 8'h80;
            20'd5535: data = 8'h80;
            20'd5536: data = 8'h7F;
            20'd5537: data = 8'h7F;
            20'd5538: data = 8'h80;
            20'd5539: data = 8'h80;
            20'd5540: data = 8'h80;
            20'd5541: data = 8'h80;
            20'd5542: data = 8'h80;
            20'd5543: data = 8'h7F;
            20'd5544: data = 8'h7F;
            20'd5545: data = 8'h80;
            20'd5546: data = 8'h7F;
            20'd5547: data = 8'h80;
            20'd5548: data = 8'h7F;
            20'd5549: data = 8'h7F;
            20'd5550: data = 8'h80;
            20'd5551: data = 8'h80;
            20'd5552: data = 8'h7F;
            20'd5553: data = 8'h7F;
            20'd5554: data = 8'h80;
            20'd5555: data = 8'h80;
            20'd5556: data = 8'h80;
            20'd5557: data = 8'h7F;
            20'd5558: data = 8'h80;
            20'd5559: data = 8'h80;
            20'd5560: data = 8'h80;
            20'd5561: data = 8'h80;
            20'd5562: data = 8'h80;
            20'd5563: data = 8'h7F;
            20'd5564: data = 8'h80;
            20'd5565: data = 8'h80;
            20'd5566: data = 8'h7F;
            20'd5567: data = 8'h80;
            20'd5568: data = 8'h80;
            20'd5569: data = 8'h7F;
            20'd5570: data = 8'h7F;
            20'd5571: data = 8'h80;
            20'd5572: data = 8'h80;
            20'd5573: data = 8'h7F;
            20'd5574: data = 8'h7F;
            20'd5575: data = 8'h80;
            20'd5576: data = 8'h80;
            20'd5577: data = 8'h7F;
            20'd5578: data = 8'h80;
            20'd5579: data = 8'h80;
            20'd5580: data = 8'h80;
            20'd5581: data = 8'h7F;
            20'd5582: data = 8'h7F;
            20'd5583: data = 8'h80;
            20'd5584: data = 8'h7F;
            20'd5585: data = 8'h80;
            20'd5586: data = 8'h80;
            20'd5587: data = 8'h7F;
            20'd5588: data = 8'h7F;
            20'd5589: data = 8'h80;
            20'd5590: data = 8'h80;
            20'd5591: data = 8'h7F;
            20'd5592: data = 8'h7F;
            20'd5593: data = 8'h7F;
            20'd5594: data = 8'h7F;
            20'd5595: data = 8'h7F;
            20'd5596: data = 8'h80;
            20'd5597: data = 8'h80;
            20'd5598: data = 8'h7F;
            20'd5599: data = 8'h80;
            20'd5600: data = 8'h7F;
            20'd5601: data = 8'h80;
            20'd5602: data = 8'h80;
            20'd5603: data = 8'h80;
            20'd5604: data = 8'h7F;
            20'd5605: data = 8'h7F;
            20'd5606: data = 8'h80;
            20'd5607: data = 8'h80;
            20'd5608: data = 8'h80;
            20'd5609: data = 8'h7F;
            20'd5610: data = 8'h7F;
            20'd5611: data = 8'h7F;
            20'd5612: data = 8'h80;
            20'd5613: data = 8'h80;
            20'd5614: data = 8'h80;
            20'd5615: data = 8'h7F;
            20'd5616: data = 8'h80;
            20'd5617: data = 8'h80;
            20'd5618: data = 8'h7F;
            20'd5619: data = 8'h7F;
            20'd5620: data = 8'h80;
            20'd5621: data = 8'h80;
            20'd5622: data = 8'h7F;
            20'd5623: data = 8'h7F;
            20'd5624: data = 8'h80;
            20'd5625: data = 8'h80;
            20'd5626: data = 8'h7F;
            20'd5627: data = 8'h80;
            20'd5628: data = 8'h80;
            20'd5629: data = 8'h80;
            20'd5630: data = 8'h7F;
            20'd5631: data = 8'h7F;
            20'd5632: data = 8'h80;
            20'd5633: data = 8'h80;
            20'd5634: data = 8'h7F;
            20'd5635: data = 8'h7F;
            20'd5636: data = 8'h80;
            20'd5637: data = 8'h7F;
            20'd5638: data = 8'h7F;
            20'd5639: data = 8'h80;
            20'd5640: data = 8'h7F;
            20'd5641: data = 8'h80;
            20'd5642: data = 8'h7F;
            20'd5643: data = 8'h80;
            20'd5644: data = 8'h7F;
            20'd5645: data = 8'h80;
            20'd5646: data = 8'h80;
            20'd5647: data = 8'h7F;
            20'd5648: data = 8'h7F;
            20'd5649: data = 8'h7F;
            20'd5650: data = 8'h7F;
            20'd5651: data = 8'h80;
            20'd5652: data = 8'h80;
            20'd5653: data = 8'h80;
            20'd5654: data = 8'h80;
            20'd5655: data = 8'h7F;
            20'd5656: data = 8'h80;
            20'd5657: data = 8'h80;
            20'd5658: data = 8'h7F;
            20'd5659: data = 8'h80;
            20'd5660: data = 8'h80;
            20'd5661: data = 8'h7F;
            20'd5662: data = 8'h80;
            20'd5663: data = 8'h80;
            20'd5664: data = 8'h7F;
            20'd5665: data = 8'h80;
            20'd5666: data = 8'h80;
            20'd5667: data = 8'h7F;
            20'd5668: data = 8'h7F;
            20'd5669: data = 8'h80;
            20'd5670: data = 8'h7F;
            20'd5671: data = 8'h80;
            20'd5672: data = 8'h7F;
            20'd5673: data = 8'h7F;
            20'd5674: data = 8'h80;
            20'd5675: data = 8'h7F;
            20'd5676: data = 8'h80;
            20'd5677: data = 8'h7F;
            20'd5678: data = 8'h80;
            20'd5679: data = 8'h7F;
            20'd5680: data = 8'h80;
            20'd5681: data = 8'h80;
            20'd5682: data = 8'h80;
            20'd5683: data = 8'h80;
            20'd5684: data = 8'h7F;
            20'd5685: data = 8'h7F;
            20'd5686: data = 8'h80;
            20'd5687: data = 8'h7F;
            20'd5688: data = 8'h80;
            20'd5689: data = 8'h7F;
            20'd5690: data = 8'h80;
            20'd5691: data = 8'h80;
            20'd5692: data = 8'h80;
            20'd5693: data = 8'h7F;
            20'd5694: data = 8'h80;
            20'd5695: data = 8'h80;
            20'd5696: data = 8'h7F;
            20'd5697: data = 8'h80;
            20'd5698: data = 8'h80;
            20'd5699: data = 8'h80;
            20'd5700: data = 8'h7F;
            20'd5701: data = 8'h7F;
            20'd5702: data = 8'h80;
            20'd5703: data = 8'h80;
            20'd5704: data = 8'h80;
            20'd5705: data = 8'h80;
            20'd5706: data = 8'h7F;
            20'd5707: data = 8'h80;
            20'd5708: data = 8'h80;
            20'd5709: data = 8'h7F;
            20'd5710: data = 8'h7F;
            20'd5711: data = 8'h80;
            20'd5712: data = 8'h80;
            20'd5713: data = 8'h80;
            20'd5714: data = 8'h80;
            20'd5715: data = 8'h7F;
            20'd5716: data = 8'h80;
            20'd5717: data = 8'h80;
            20'd5718: data = 8'h7F;
            20'd5719: data = 8'h80;
            20'd5720: data = 8'h80;
            20'd5721: data = 8'h7F;
            20'd5722: data = 8'h7F;
            20'd5723: data = 8'h80;
            20'd5724: data = 8'h80;
            20'd5725: data = 8'h80;
            20'd5726: data = 8'h7F;
            20'd5727: data = 8'h80;
            20'd5728: data = 8'h80;
            20'd5729: data = 8'h80;
            20'd5730: data = 8'h80;
            20'd5731: data = 8'h80;
            20'd5732: data = 8'h7F;
            20'd5733: data = 8'h80;
            20'd5734: data = 8'h80;
            20'd5735: data = 8'h80;
            20'd5736: data = 8'h7F;
            20'd5737: data = 8'h80;
            20'd5738: data = 8'h7F;
            20'd5739: data = 8'h80;
            20'd5740: data = 8'h80;
            20'd5741: data = 8'h80;
            20'd5742: data = 8'h7F;
            20'd5743: data = 8'h80;
            20'd5744: data = 8'h80;
            20'd5745: data = 8'h80;
            20'd5746: data = 8'h80;
            20'd5747: data = 8'h80;
            20'd5748: data = 8'h80;
            20'd5749: data = 8'h80;
            20'd5750: data = 8'h7F;
            20'd5751: data = 8'h80;
            20'd5752: data = 8'h7F;
            20'd5753: data = 8'h80;
            20'd5754: data = 8'h80;
            20'd5755: data = 8'h7F;
            20'd5756: data = 8'h80;
            20'd5757: data = 8'h7F;
            20'd5758: data = 8'h7F;
            20'd5759: data = 8'h80;
            20'd5760: data = 8'h80;
            20'd5761: data = 8'h80;
            20'd5762: data = 8'h80;
            20'd5763: data = 8'h80;
            20'd5764: data = 8'h7F;
            20'd5765: data = 8'h7F;
            20'd5766: data = 8'h80;
            20'd5767: data = 8'h80;
            20'd5768: data = 8'h80;
            20'd5769: data = 8'h80;
            20'd5770: data = 8'h7F;
            20'd5771: data = 8'h80;
            20'd5772: data = 8'h80;
            20'd5773: data = 8'h80;
            20'd5774: data = 8'h80;
            20'd5775: data = 8'h80;
            20'd5776: data = 8'h80;
            20'd5777: data = 8'h80;
            20'd5778: data = 8'h80;
            20'd5779: data = 8'h80;
            20'd5780: data = 8'h80;
            20'd5781: data = 8'h80;
            20'd5782: data = 8'h7F;
            20'd5783: data = 8'h7F;
            20'd5784: data = 8'h80;
            20'd5785: data = 8'h80;
            20'd5786: data = 8'h80;
            20'd5787: data = 8'h7F;
            20'd5788: data = 8'h80;
            20'd5789: data = 8'h7F;
            20'd5790: data = 8'h7F;
            20'd5791: data = 8'h80;
            20'd5792: data = 8'h80;
            20'd5793: data = 8'h80;
            20'd5794: data = 8'h80;
            20'd5795: data = 8'h7F;
            20'd5796: data = 8'h80;
            20'd5797: data = 8'h7F;
            20'd5798: data = 8'h80;
            20'd5799: data = 8'h80;
            20'd5800: data = 8'h80;
            20'd5801: data = 8'h7F;
            20'd5802: data = 8'h7F;
            20'd5803: data = 8'h80;
            20'd5804: data = 8'h80;
            20'd5805: data = 8'h7F;
            20'd5806: data = 8'h80;
            20'd5807: data = 8'h80;
            20'd5808: data = 8'h80;
            20'd5809: data = 8'h80;
            20'd5810: data = 8'h80;
            20'd5811: data = 8'h80;
            20'd5812: data = 8'h80;
            20'd5813: data = 8'h80;
            20'd5814: data = 8'h7F;
            20'd5815: data = 8'h80;
            20'd5816: data = 8'h80;
            20'd5817: data = 8'h80;
            20'd5818: data = 8'h80;
            20'd5819: data = 8'h80;
            20'd5820: data = 8'h7F;
            20'd5821: data = 8'h80;
            20'd5822: data = 8'h7F;
            20'd5823: data = 8'h80;
            20'd5824: data = 8'h80;
            20'd5825: data = 8'h80;
            20'd5826: data = 8'h7F;
            20'd5827: data = 8'h80;
            20'd5828: data = 8'h7F;
            20'd5829: data = 8'h80;
            20'd5830: data = 8'h80;
            20'd5831: data = 8'h80;
            20'd5832: data = 8'h80;
            20'd5833: data = 8'h80;
            20'd5834: data = 8'h80;
            20'd5835: data = 8'h80;
            20'd5836: data = 8'h80;
            20'd5837: data = 8'h7F;
            20'd5838: data = 8'h80;
            20'd5839: data = 8'h80;
            20'd5840: data = 8'h80;
            20'd5841: data = 8'h80;
            20'd5842: data = 8'h7F;
            20'd5843: data = 8'h80;
            20'd5844: data = 8'h80;
            20'd5845: data = 8'h80;
            20'd5846: data = 8'h80;
            20'd5847: data = 8'h80;
            20'd5848: data = 8'h80;
            20'd5849: data = 8'h7F;
            20'd5850: data = 8'h80;
            20'd5851: data = 8'h80;
            20'd5852: data = 8'h80;
            20'd5853: data = 8'h80;
            20'd5854: data = 8'h80;
            20'd5855: data = 8'h80;
            20'd5856: data = 8'h80;
            20'd5857: data = 8'h80;
            20'd5858: data = 8'h80;
            20'd5859: data = 8'h80;
            20'd5860: data = 8'h80;
            20'd5861: data = 8'h80;
            20'd5862: data = 8'h80;
            20'd5863: data = 8'h80;
            20'd5864: data = 8'h80;
            20'd5865: data = 8'h80;
            20'd5866: data = 8'h80;
            20'd5867: data = 8'h80;
            20'd5868: data = 8'h80;
            20'd5869: data = 8'h80;
            20'd5870: data = 8'h7F;
            20'd5871: data = 8'h80;
            20'd5872: data = 8'h80;
            20'd5873: data = 8'h80;
            20'd5874: data = 8'h7F;
            20'd5875: data = 8'h80;
            20'd5876: data = 8'h80;
            20'd5877: data = 8'h80;
            20'd5878: data = 8'h80;
            20'd5879: data = 8'h80;
            20'd5880: data = 8'h80;
            20'd5881: data = 8'h80;
            20'd5882: data = 8'h80;
            20'd5883: data = 8'h7F;
            20'd5884: data = 8'h80;
            20'd5885: data = 8'h80;
            20'd5886: data = 8'h80;
            20'd5887: data = 8'h80;
            20'd5888: data = 8'h80;
            20'd5889: data = 8'h80;
            20'd5890: data = 8'h80;
            20'd5891: data = 8'h80;
            20'd5892: data = 8'h80;
            20'd5893: data = 8'h80;
            20'd5894: data = 8'h80;
            20'd5895: data = 8'h80;
            20'd5896: data = 8'h80;
            20'd5897: data = 8'h80;
            20'd5898: data = 8'h80;
            20'd5899: data = 8'h80;
            20'd5900: data = 8'h80;
            20'd5901: data = 8'h80;
            20'd5902: data = 8'h80;
            20'd5903: data = 8'h80;
            20'd5904: data = 8'h80;
            20'd5905: data = 8'h80;
            20'd5906: data = 8'h80;
            20'd5907: data = 8'h80;
            20'd5908: data = 8'h80;
            20'd5909: data = 8'h80;
            20'd5910: data = 8'h80;
            20'd5911: data = 8'h80;
            20'd5912: data = 8'h80;
            20'd5913: data = 8'h80;
            20'd5914: data = 8'h80;
            20'd5915: data = 8'h80;
            20'd5916: data = 8'h80;
            20'd5917: data = 8'h80;
            20'd5918: data = 8'h80;
            20'd5919: data = 8'h80;
            20'd5920: data = 8'h80;
            20'd5921: data = 8'h7F;
            20'd5922: data = 8'h80;
            20'd5923: data = 8'h80;
            20'd5924: data = 8'h80;
            20'd5925: data = 8'h80;
            20'd5926: data = 8'h80;
            20'd5927: data = 8'h80;
            20'd5928: data = 8'h80;
            20'd5929: data = 8'h80;
            20'd5930: data = 8'h80;
            20'd5931: data = 8'h80;
            20'd5932: data = 8'h80;
            20'd5933: data = 8'h80;
            20'd5934: data = 8'h80;
            20'd5935: data = 8'h80;
            20'd5936: data = 8'h80;
            20'd5937: data = 8'h80;
            20'd5938: data = 8'h80;
            20'd5939: data = 8'h80;
            20'd5940: data = 8'h80;
            20'd5941: data = 8'h80;
            20'd5942: data = 8'h80;
            20'd5943: data = 8'h80;
            20'd5944: data = 8'h80;
            20'd5945: data = 8'h80;
            20'd5946: data = 8'h80;
            20'd5947: data = 8'h80;
            20'd5948: data = 8'h80;
            20'd5949: data = 8'h80;
            20'd5950: data = 8'h80;
            20'd5951: data = 8'h80;
            20'd5952: data = 8'h80;
            20'd5953: data = 8'h80;
            20'd5954: data = 8'h80;
            20'd5955: data = 8'h80;
            20'd5956: data = 8'h80;
            20'd5957: data = 8'h80;
            20'd5958: data = 8'h80;
            20'd5959: data = 8'h80;
            20'd5960: data = 8'h80;
            20'd5961: data = 8'h80;
            20'd5962: data = 8'h80;
            20'd5963: data = 8'h80;
            20'd5964: data = 8'h80;
            20'd5965: data = 8'h80;
            20'd5966: data = 8'h80;
            20'd5967: data = 8'h80;
            20'd5968: data = 8'h80;
            20'd5969: data = 8'h80;
            20'd5970: data = 8'h80;
            20'd5971: data = 8'h80;
            20'd5972: data = 8'h80;
            20'd5973: data = 8'h80;
            20'd5974: data = 8'h80;
            20'd5975: data = 8'h80;
            20'd5976: data = 8'h80;
            20'd5977: data = 8'h80;
            20'd5978: data = 8'h80;
            20'd5979: data = 8'h80;
            20'd5980: data = 8'h80;
            20'd5981: data = 8'h80;
            20'd5982: data = 8'h80;
            20'd5983: data = 8'h80;
            20'd5984: data = 8'h80;
            20'd5985: data = 8'h80;
            20'd5986: data = 8'h80;
            20'd5987: data = 8'h80;
            20'd5988: data = 8'h80;
            20'd5989: data = 8'h80;
            20'd5990: data = 8'h80;
            20'd5991: data = 8'h80;
            20'd5992: data = 8'h80;
            20'd5993: data = 8'h80;
            20'd5994: data = 8'h80;
            20'd5995: data = 8'h80;
            20'd5996: data = 8'h80;
            20'd5997: data = 8'h80;
            20'd5998: data = 8'h80;
            20'd5999: data = 8'h80;
            20'd6000: data = 8'h80;
            20'd6001: data = 8'h80;
            20'd6002: data = 8'h80;
            20'd6003: data = 8'h80;
            20'd6004: data = 8'h80;
            20'd6005: data = 8'h80;
            20'd6006: data = 8'h80;
            20'd6007: data = 8'h80;
            20'd6008: data = 8'h80;
            20'd6009: data = 8'h80;
            20'd6010: data = 8'h80;
            20'd6011: data = 8'h80;
            20'd6012: data = 8'h80;
            20'd6013: data = 8'h80;
            20'd6014: data = 8'h80;
            20'd6015: data = 8'h80;
            20'd6016: data = 8'h80;
            20'd6017: data = 8'h80;
            20'd6018: data = 8'h80;
            20'd6019: data = 8'h80;
            20'd6020: data = 8'h80;
            20'd6021: data = 8'h80;
            20'd6022: data = 8'h80;
            20'd6023: data = 8'h80;
            20'd6024: data = 8'h80;
            20'd6025: data = 8'h80;
            20'd6026: data = 8'h80;
            20'd6027: data = 8'h80;
            20'd6028: data = 8'h80;
            20'd6029: data = 8'h80;
            20'd6030: data = 8'h80;
            20'd6031: data = 8'h80;
            20'd6032: data = 8'h80;
            20'd6033: data = 8'h80;
            20'd6034: data = 8'h80;
            20'd6035: data = 8'h80;
            20'd6036: data = 8'h80;
            20'd6037: data = 8'h80;
            20'd6038: data = 8'h80;
            20'd6039: data = 8'h80;
            20'd6040: data = 8'h80;
            20'd6041: data = 8'h80;
            20'd6042: data = 8'h80;
            20'd6043: data = 8'h80;
            20'd6044: data = 8'h80;
            20'd6045: data = 8'h80;
            20'd6046: data = 8'h80;
            20'd6047: data = 8'h80;
            20'd6048: data = 8'h80;
            20'd6049: data = 8'h80;
            20'd6050: data = 8'h80;
            20'd6051: data = 8'h80;
            20'd6052: data = 8'h80;
            20'd6053: data = 8'h80;
            20'd6054: data = 8'h80;
            20'd6055: data = 8'h80;
            20'd6056: data = 8'h80;
            20'd6057: data = 8'h80;
            20'd6058: data = 8'h80;
            20'd6059: data = 8'h80;
            20'd6060: data = 8'h80;
            20'd6061: data = 8'h80;
            20'd6062: data = 8'h80;
            20'd6063: data = 8'h80;
            20'd6064: data = 8'h80;
            20'd6065: data = 8'h80;
            20'd6066: data = 8'h80;
            20'd6067: data = 8'h80;
            20'd6068: data = 8'h80;
            20'd6069: data = 8'h80;
            20'd6070: data = 8'h80;
            20'd6071: data = 8'h80;
            20'd6072: data = 8'h80;
            20'd6073: data = 8'h80;
            20'd6074: data = 8'h80;
            20'd6075: data = 8'h80;
            20'd6076: data = 8'h80;
            20'd6077: data = 8'h80;
            20'd6078: data = 8'h80;
            20'd6079: data = 8'h80;
            20'd6080: data = 8'h80;
            20'd6081: data = 8'h80;
            20'd6082: data = 8'h80;
            20'd6083: data = 8'h80;
            20'd6084: data = 8'h80;
            20'd6085: data = 8'h80;
            20'd6086: data = 8'h80;
            20'd6087: data = 8'h80;
            20'd6088: data = 8'h80;
            20'd6089: data = 8'h80;
            20'd6090: data = 8'h80;
            20'd6091: data = 8'h80;
            20'd6092: data = 8'h80;
            20'd6093: data = 8'h80;
            20'd6094: data = 8'h80;
            20'd6095: data = 8'h80;
            20'd6096: data = 8'h80;
            20'd6097: data = 8'h80;
            20'd6098: data = 8'h80;
            20'd6099: data = 8'h80;
            20'd6100: data = 8'h80;
            20'd6101: data = 8'h80;
            20'd6102: data = 8'h80;
            20'd6103: data = 8'h80;
            20'd6104: data = 8'h80;
            20'd6105: data = 8'h80;
            20'd6106: data = 8'h80;
            20'd6107: data = 8'h80;
            20'd6108: data = 8'h80;
            20'd6109: data = 8'h80;
            20'd6110: data = 8'h80;
            20'd6111: data = 8'h80;
            20'd6112: data = 8'h80;
            20'd6113: data = 8'h80;
            20'd6114: data = 8'h80;
            20'd6115: data = 8'h80;
            20'd6116: data = 8'h80;
            20'd6117: data = 8'h80;
            20'd6118: data = 8'h80;
            20'd6119: data = 8'h80;
            20'd6120: data = 8'h80;
            20'd6121: data = 8'h80;
            20'd6122: data = 8'h80;
            20'd6123: data = 8'h80;
            20'd6124: data = 8'h80;
            20'd6125: data = 8'h80;
            20'd6126: data = 8'h80;
            20'd6127: data = 8'h80;
            20'd6128: data = 8'h80;
            20'd6129: data = 8'h80;
            20'd6130: data = 8'h80;
            20'd6131: data = 8'h80;
            20'd6132: data = 8'h80;
            20'd6133: data = 8'h80;
            20'd6134: data = 8'h80;
            20'd6135: data = 8'h80;
            20'd6136: data = 8'h80;
            20'd6137: data = 8'h80;
            20'd6138: data = 8'h80;
            20'd6139: data = 8'h80;
            20'd6140: data = 8'h80;
            20'd6141: data = 8'h80;
            20'd6142: data = 8'h80;
            20'd6143: data = 8'h80;
            20'd6144: data = 8'h80;
            20'd6145: data = 8'h80;
            20'd6146: data = 8'h80;
            20'd6147: data = 8'h80;
            20'd6148: data = 8'h80;
            20'd6149: data = 8'h80;
            20'd6150: data = 8'h80;
            20'd6151: data = 8'h80;
            20'd6152: data = 8'h80;
            20'd6153: data = 8'h80;
            20'd6154: data = 8'h80;
            20'd6155: data = 8'h80;
            20'd6156: data = 8'h80;
            20'd6157: data = 8'h80;
            20'd6158: data = 8'h80;
            20'd6159: data = 8'h80;
            20'd6160: data = 8'h80;
            20'd6161: data = 8'h80;
            20'd6162: data = 8'h80;
            20'd6163: data = 8'h80;
            20'd6164: data = 8'h80;
            20'd6165: data = 8'h80;
            20'd6166: data = 8'h80;
            20'd6167: data = 8'h80;
            20'd6168: data = 8'h80;
            20'd6169: data = 8'h80;
            20'd6170: data = 8'h80;
            20'd6171: data = 8'h80;
            20'd6172: data = 8'h80;
            20'd6173: data = 8'h80;
            20'd6174: data = 8'h80;
            20'd6175: data = 8'h80;
            20'd6176: data = 8'h80;
            20'd6177: data = 8'h80;
            20'd6178: data = 8'h80;
            20'd6179: data = 8'h80;
            20'd6180: data = 8'h80;
            20'd6181: data = 8'h80;
            20'd6182: data = 8'h80;
            20'd6183: data = 8'h80;
            20'd6184: data = 8'h80;
            20'd6185: data = 8'h80;
            20'd6186: data = 8'h80;
            20'd6187: data = 8'h80;
            20'd6188: data = 8'h80;
            20'd6189: data = 8'h80;
            20'd6190: data = 8'h80;
            20'd6191: data = 8'h80;
            20'd6192: data = 8'h80;
            20'd6193: data = 8'h80;
            20'd6194: data = 8'h80;
            20'd6195: data = 8'h80;
            20'd6196: data = 8'h80;
            20'd6197: data = 8'h80;
            20'd6198: data = 8'h80;
            20'd6199: data = 8'h80;
            20'd6200: data = 8'h80;
            20'd6201: data = 8'h80;
            20'd6202: data = 8'h80;
            20'd6203: data = 8'h80;
            20'd6204: data = 8'h80;
            20'd6205: data = 8'h80;
            20'd6206: data = 8'h80;
            20'd6207: data = 8'h80;
            20'd6208: data = 8'h80;
            20'd6209: data = 8'h80;
            20'd6210: data = 8'h80;
            20'd6211: data = 8'h80;
            20'd6212: data = 8'h80;
            20'd6213: data = 8'h80;
            20'd6214: data = 8'h80;
            20'd6215: data = 8'h80;
            20'd6216: data = 8'h80;
            20'd6217: data = 8'h80;
            20'd6218: data = 8'h80;
            20'd6219: data = 8'h80;
            20'd6220: data = 8'h80;
            20'd6221: data = 8'h80;
            20'd6222: data = 8'h80;
            20'd6223: data = 8'h80;
            20'd6224: data = 8'h80;
            20'd6225: data = 8'h80;
            20'd6226: data = 8'h80;
            20'd6227: data = 8'h80;
            20'd6228: data = 8'h80;
            20'd6229: data = 8'h80;
            20'd6230: data = 8'h80;
            20'd6231: data = 8'h80;
            20'd6232: data = 8'h80;
            20'd6233: data = 8'h80;
            20'd6234: data = 8'h80;
            20'd6235: data = 8'h80;
            20'd6236: data = 8'h80;
            20'd6237: data = 8'h80;
            20'd6238: data = 8'h80;
            20'd6239: data = 8'h80;
            20'd6240: data = 8'h80;
            20'd6241: data = 8'h80;
            20'd6242: data = 8'h80;
            20'd6243: data = 8'h80;
            20'd6244: data = 8'h80;
            20'd6245: data = 8'h80;
            20'd6246: data = 8'h80;
            20'd6247: data = 8'h80;
            20'd6248: data = 8'h80;
            20'd6249: data = 8'h80;
            20'd6250: data = 8'h80;
            20'd6251: data = 8'h80;
            20'd6252: data = 8'h80;
            20'd6253: data = 8'h80;
            20'd6254: data = 8'h80;
            20'd6255: data = 8'h80;
            20'd6256: data = 8'h80;
            20'd6257: data = 8'h80;
            20'd6258: data = 8'h80;
            20'd6259: data = 8'h80;
            20'd6260: data = 8'h80;
            20'd6261: data = 8'h80;
            20'd6262: data = 8'h80;
            20'd6263: data = 8'h80;
            20'd6264: data = 8'h80;
            20'd6265: data = 8'h80;
            20'd6266: data = 8'h80;
            20'd6267: data = 8'h80;
            20'd6268: data = 8'h80;
            20'd6269: data = 8'h80;
            20'd6270: data = 8'h80;
            20'd6271: data = 8'h80;
            20'd6272: data = 8'h80;
            20'd6273: data = 8'h80;
            20'd6274: data = 8'h80;
            20'd6275: data = 8'h80;
            20'd6276: data = 8'h80;
            20'd6277: data = 8'h80;
            20'd6278: data = 8'h80;
            20'd6279: data = 8'h80;
            20'd6280: data = 8'h80;
            20'd6281: data = 8'h80;
            20'd6282: data = 8'h80;
            20'd6283: data = 8'h80;
            20'd6284: data = 8'h80;
            20'd6285: data = 8'h80;
            20'd6286: data = 8'h80;
            20'd6287: data = 8'h80;
            20'd6288: data = 8'h80;
            20'd6289: data = 8'h80;
            20'd6290: data = 8'h80;
            20'd6291: data = 8'h80;
            20'd6292: data = 8'h80;
            20'd6293: data = 8'h80;
            20'd6294: data = 8'h80;
            20'd6295: data = 8'h80;
            20'd6296: data = 8'h80;
            20'd6297: data = 8'h80;
            20'd6298: data = 8'h80;
            20'd6299: data = 8'h80;
            20'd6300: data = 8'h80;
            20'd6301: data = 8'h80;
            20'd6302: data = 8'h80;
            20'd6303: data = 8'h80;
            20'd6304: data = 8'h80;
            20'd6305: data = 8'h80;
            20'd6306: data = 8'h80;
            20'd6307: data = 8'h80;
            20'd6308: data = 8'h80;
            20'd6309: data = 8'h80;
            20'd6310: data = 8'h80;
            20'd6311: data = 8'h80;
            20'd6312: data = 8'h80;
            20'd6313: data = 8'h80;
            20'd6314: data = 8'h80;
            20'd6315: data = 8'h80;
            20'd6316: data = 8'h80;
            20'd6317: data = 8'h80;
            20'd6318: data = 8'h80;
            20'd6319: data = 8'h80;
            20'd6320: data = 8'h80;
            20'd6321: data = 8'h80;
            20'd6322: data = 8'h80;
            20'd6323: data = 8'h80;
            20'd6324: data = 8'h80;
            20'd6325: data = 8'h80;
            20'd6326: data = 8'h80;
            20'd6327: data = 8'h80;
            20'd6328: data = 8'h80;
            20'd6329: data = 8'h80;
            20'd6330: data = 8'h80;
            20'd6331: data = 8'h80;
            20'd6332: data = 8'h80;
            20'd6333: data = 8'h80;
            20'd6334: data = 8'h80;
            20'd6335: data = 8'h80;
            20'd6336: data = 8'h80;
            20'd6337: data = 8'h80;
            20'd6338: data = 8'h80;
            20'd6339: data = 8'h80;
            20'd6340: data = 8'h80;
            20'd6341: data = 8'h80;
            20'd6342: data = 8'h80;
            20'd6343: data = 8'h80;
            20'd6344: data = 8'h80;
            20'd6345: data = 8'h80;
            20'd6346: data = 8'h80;
            20'd6347: data = 8'h80;
            20'd6348: data = 8'h80;
            20'd6349: data = 8'h80;
            20'd6350: data = 8'h80;
            20'd6351: data = 8'h80;
            20'd6352: data = 8'h80;
            20'd6353: data = 8'h80;
            20'd6354: data = 8'h80;
            20'd6355: data = 8'h80;
            20'd6356: data = 8'h80;
            20'd6357: data = 8'h80;
            20'd6358: data = 8'h80;
            20'd6359: data = 8'h80;
            20'd6360: data = 8'h80;
            20'd6361: data = 8'h80;
            20'd6362: data = 8'h80;
            20'd6363: data = 8'h80;
            20'd6364: data = 8'h80;
            20'd6365: data = 8'h80;
            20'd6366: data = 8'h80;
            20'd6367: data = 8'h80;
            20'd6368: data = 8'h80;
            20'd6369: data = 8'h80;
            20'd6370: data = 8'h80;
            20'd6371: data = 8'h80;
            20'd6372: data = 8'h80;
            20'd6373: data = 8'h80;
            20'd6374: data = 8'h80;
            20'd6375: data = 8'h80;
            20'd6376: data = 8'h80;
            20'd6377: data = 8'h80;
            20'd6378: data = 8'h80;
            20'd6379: data = 8'h80;
            20'd6380: data = 8'h80;
            20'd6381: data = 8'h80;
            20'd6382: data = 8'h80;
            20'd6383: data = 8'h80;
            20'd6384: data = 8'h80;
            20'd6385: data = 8'h80;
            20'd6386: data = 8'h80;
            20'd6387: data = 8'h80;
            20'd6388: data = 8'h80;
            20'd6389: data = 8'h80;
            20'd6390: data = 8'h80;
            20'd6391: data = 8'h80;
            20'd6392: data = 8'h80;
            20'd6393: data = 8'h80;
            20'd6394: data = 8'h80;
            20'd6395: data = 8'h80;
            20'd6396: data = 8'h80;
            20'd6397: data = 8'h80;
            20'd6398: data = 8'h80;
            20'd6399: data = 8'h80;
            20'd6400: data = 8'h80;
            20'd6401: data = 8'h80;
            20'd6402: data = 8'h80;
            20'd6403: data = 8'h80;
            20'd6404: data = 8'h80;
            20'd6405: data = 8'h80;
            20'd6406: data = 8'h80;
            20'd6407: data = 8'h80;
            20'd6408: data = 8'h80;
            20'd6409: data = 8'h80;
            20'd6410: data = 8'h80;
            20'd6411: data = 8'h80;
            20'd6412: data = 8'h80;
            20'd6413: data = 8'h80;
            20'd6414: data = 8'h80;
            20'd6415: data = 8'h80;
            20'd6416: data = 8'h80;
            20'd6417: data = 8'h80;
            20'd6418: data = 8'h80;
            20'd6419: data = 8'h80;
            20'd6420: data = 8'h80;
            20'd6421: data = 8'h80;
            20'd6422: data = 8'h80;
            20'd6423: data = 8'h80;
            20'd6424: data = 8'h80;
            20'd6425: data = 8'h80;
            20'd6426: data = 8'h80;
            20'd6427: data = 8'h80;
            20'd6428: data = 8'h80;
            20'd6429: data = 8'h80;
            20'd6430: data = 8'h80;
            20'd6431: data = 8'h80;
            20'd6432: data = 8'h80;
            20'd6433: data = 8'h80;
            20'd6434: data = 8'h80;
            20'd6435: data = 8'h80;
            20'd6436: data = 8'h80;
            20'd6437: data = 8'h80;
            20'd6438: data = 8'h80;
            20'd6439: data = 8'h80;
            20'd6440: data = 8'h80;
            20'd6441: data = 8'h80;
            20'd6442: data = 8'h80;
            20'd6443: data = 8'h80;
            20'd6444: data = 8'h80;
            20'd6445: data = 8'h80;
            20'd6446: data = 8'h80;
            20'd6447: data = 8'h80;
            20'd6448: data = 8'h80;
            20'd6449: data = 8'h80;
            20'd6450: data = 8'h80;
            20'd6451: data = 8'h80;
            20'd6452: data = 8'h80;
            20'd6453: data = 8'h80;
            20'd6454: data = 8'h80;
            20'd6455: data = 8'h80;
            20'd6456: data = 8'h80;
            20'd6457: data = 8'h80;
            20'd6458: data = 8'h80;
            20'd6459: data = 8'h80;
            20'd6460: data = 8'h80;
            20'd6461: data = 8'h80;
            20'd6462: data = 8'h80;
            20'd6463: data = 8'h80;
            20'd6464: data = 8'h80;
            20'd6465: data = 8'h80;
            20'd6466: data = 8'h80;
            20'd6467: data = 8'h80;
            20'd6468: data = 8'h80;
            20'd6469: data = 8'h80;
            20'd6470: data = 8'h80;
            20'd6471: data = 8'h80;
            20'd6472: data = 8'h80;
            20'd6473: data = 8'h80;
            20'd6474: data = 8'h80;
            20'd6475: data = 8'h80;
            20'd6476: data = 8'h80;
            20'd6477: data = 8'h80;
            20'd6478: data = 8'h80;
            20'd6479: data = 8'h80;
            20'd6480: data = 8'h80;
            20'd6481: data = 8'h80;
            20'd6482: data = 8'h80;
            20'd6483: data = 8'h80;
            20'd6484: data = 8'h80;
            20'd6485: data = 8'h80;
            20'd6486: data = 8'h80;
            20'd6487: data = 8'h80;
            20'd6488: data = 8'h80;
            20'd6489: data = 8'h80;
            20'd6490: data = 8'h80;
            20'd6491: data = 8'h80;
            20'd6492: data = 8'h80;
            20'd6493: data = 8'h80;
            20'd6494: data = 8'h80;
            20'd6495: data = 8'h80;
            20'd6496: data = 8'h80;
            20'd6497: data = 8'h80;
            20'd6498: data = 8'h80;
            20'd6499: data = 8'h80;
            20'd6500: data = 8'h80;
            20'd6501: data = 8'h80;
            20'd6502: data = 8'h80;
            20'd6503: data = 8'h80;
            20'd6504: data = 8'h80;
            20'd6505: data = 8'h80;
            20'd6506: data = 8'h80;
            20'd6507: data = 8'h80;
            20'd6508: data = 8'h80;
            20'd6509: data = 8'h80;
            20'd6510: data = 8'h80;
            20'd6511: data = 8'h80;
            20'd6512: data = 8'h80;
            20'd6513: data = 8'h80;
            20'd6514: data = 8'h80;
            20'd6515: data = 8'h80;
            20'd6516: data = 8'h80;
            20'd6517: data = 8'h80;
            20'd6518: data = 8'h80;
            20'd6519: data = 8'h80;
            20'd6520: data = 8'h80;
            20'd6521: data = 8'h80;
            20'd6522: data = 8'h80;
            20'd6523: data = 8'h80;
            20'd6524: data = 8'h80;
            20'd6525: data = 8'h80;
            20'd6526: data = 8'h80;
            20'd6527: data = 8'h80;
            20'd6528: data = 8'h80;
            20'd6529: data = 8'h80;
            20'd6530: data = 8'h80;
            20'd6531: data = 8'h80;
            20'd6532: data = 8'h80;
            20'd6533: data = 8'h80;
            20'd6534: data = 8'h80;
            20'd6535: data = 8'h80;
            20'd6536: data = 8'h80;
            20'd6537: data = 8'h80;
            20'd6538: data = 8'h80;
            20'd6539: data = 8'h80;
            20'd6540: data = 8'h80;
            20'd6541: data = 8'h80;
            20'd6542: data = 8'h80;
            20'd6543: data = 8'h80;
            20'd6544: data = 8'h80;
            20'd6545: data = 8'h80;
            20'd6546: data = 8'h80;
            20'd6547: data = 8'h80;
            20'd6548: data = 8'h80;
            20'd6549: data = 8'h80;
            20'd6550: data = 8'h80;
            20'd6551: data = 8'h80;
            20'd6552: data = 8'h80;
            20'd6553: data = 8'h80;
            20'd6554: data = 8'h80;
            20'd6555: data = 8'h80;
            20'd6556: data = 8'h80;
            20'd6557: data = 8'h80;
            20'd6558: data = 8'h80;
            20'd6559: data = 8'h80;
            20'd6560: data = 8'h80;
            20'd6561: data = 8'h80;
            20'd6562: data = 8'h80;
            20'd6563: data = 8'h80;
            20'd6564: data = 8'h80;
            20'd6565: data = 8'h80;
            20'd6566: data = 8'h80;
            20'd6567: data = 8'h80;
            20'd6568: data = 8'h80;
            20'd6569: data = 8'h80;
            20'd6570: data = 8'h80;
            20'd6571: data = 8'h80;
            20'd6572: data = 8'h80;
            20'd6573: data = 8'h80;
            20'd6574: data = 8'h80;
            20'd6575: data = 8'h80;
            20'd6576: data = 8'h80;
            20'd6577: data = 8'h80;
            20'd6578: data = 8'h80;
            20'd6579: data = 8'h80;
            20'd6580: data = 8'h80;
            20'd6581: data = 8'h80;
            20'd6582: data = 8'h80;
            20'd6583: data = 8'h80;
            20'd6584: data = 8'h80;
            20'd6585: data = 8'h80;
            20'd6586: data = 8'h80;
            20'd6587: data = 8'h80;
            20'd6588: data = 8'h80;
            20'd6589: data = 8'h80;
            20'd6590: data = 8'h80;
            20'd6591: data = 8'h80;
            20'd6592: data = 8'h80;
            20'd6593: data = 8'h80;
            20'd6594: data = 8'h80;
            20'd6595: data = 8'h80;
            20'd6596: data = 8'h80;
            20'd6597: data = 8'h80;
            20'd6598: data = 8'h80;
            20'd6599: data = 8'h80;
            20'd6600: data = 8'h80;
            20'd6601: data = 8'h80;
            20'd6602: data = 8'h80;
            20'd6603: data = 8'h80;
            20'd6604: data = 8'h80;
            20'd6605: data = 8'h80;
            20'd6606: data = 8'h80;
            20'd6607: data = 8'h80;
            20'd6608: data = 8'h80;
            20'd6609: data = 8'h80;
            20'd6610: data = 8'h80;
            20'd6611: data = 8'h80;
            20'd6612: data = 8'h80;
            20'd6613: data = 8'h80;
            20'd6614: data = 8'h80;
            20'd6615: data = 8'h80;
            20'd6616: data = 8'h80;
            20'd6617: data = 8'h80;
            20'd6618: data = 8'h80;
            20'd6619: data = 8'h80;
            20'd6620: data = 8'h80;
            20'd6621: data = 8'h80;
            20'd6622: data = 8'h80;
            20'd6623: data = 8'h80;
            20'd6624: data = 8'h80;
            20'd6625: data = 8'h80;
            20'd6626: data = 8'h80;
            20'd6627: data = 8'h80;
            20'd6628: data = 8'h80;
            20'd6629: data = 8'h80;
            20'd6630: data = 8'h80;
            20'd6631: data = 8'h80;
            20'd6632: data = 8'h80;
            20'd6633: data = 8'h80;
            20'd6634: data = 8'h80;
            20'd6635: data = 8'h80;
            20'd6636: data = 8'h80;
            20'd6637: data = 8'h80;
            20'd6638: data = 8'h80;
            20'd6639: data = 8'h80;
            20'd6640: data = 8'h80;
            20'd6641: data = 8'h80;
            20'd6642: data = 8'h80;
            20'd6643: data = 8'h80;
            20'd6644: data = 8'h80;
            20'd6645: data = 8'h80;
            20'd6646: data = 8'h80;
            20'd6647: data = 8'h80;
            20'd6648: data = 8'h80;
            20'd6649: data = 8'h80;
            20'd6650: data = 8'h80;
            20'd6651: data = 8'h80;
            20'd6652: data = 8'h80;
            20'd6653: data = 8'h80;
            20'd6654: data = 8'h80;
            20'd6655: data = 8'h80;
            20'd6656: data = 8'h80;
            20'd6657: data = 8'h80;
            20'd6658: data = 8'h80;
            20'd6659: data = 8'h80;
            20'd6660: data = 8'h80;
            20'd6661: data = 8'h80;
            20'd6662: data = 8'h80;
            20'd6663: data = 8'h80;
            20'd6664: data = 8'h80;
            20'd6665: data = 8'h80;
            20'd6666: data = 8'h80;
            20'd6667: data = 8'h80;
            20'd6668: data = 8'h80;
            20'd6669: data = 8'h80;
            20'd6670: data = 8'h80;
            20'd6671: data = 8'h80;
            20'd6672: data = 8'h80;
            20'd6673: data = 8'h80;
            20'd6674: data = 8'h80;
            20'd6675: data = 8'h80;
            20'd6676: data = 8'h80;
            20'd6677: data = 8'h80;
            20'd6678: data = 8'h80;
            20'd6679: data = 8'h80;
            20'd6680: data = 8'h80;
            20'd6681: data = 8'h80;
            20'd6682: data = 8'h80;
            20'd6683: data = 8'h80;
            20'd6684: data = 8'h80;
            20'd6685: data = 8'h80;
            20'd6686: data = 8'h80;
            20'd6687: data = 8'h80;
            20'd6688: data = 8'h80;
            20'd6689: data = 8'h80;
            20'd6690: data = 8'h80;
            20'd6691: data = 8'h80;
            20'd6692: data = 8'h80;
            20'd6693: data = 8'h80;
            20'd6694: data = 8'h80;
            20'd6695: data = 8'h80;
            20'd6696: data = 8'h80;
            20'd6697: data = 8'h80;
            20'd6698: data = 8'h80;
            20'd6699: data = 8'h80;
            20'd6700: data = 8'h80;
            20'd6701: data = 8'h80;
            20'd6702: data = 8'h80;
            20'd6703: data = 8'h80;
            20'd6704: data = 8'h80;
            20'd6705: data = 8'h80;
            20'd6706: data = 8'h80;
            20'd6707: data = 8'h80;
            20'd6708: data = 8'h80;
            20'd6709: data = 8'h80;
            20'd6710: data = 8'h80;
            20'd6711: data = 8'h80;
            20'd6712: data = 8'h80;
            20'd6713: data = 8'h80;
            20'd6714: data = 8'h80;
            20'd6715: data = 8'h80;
            20'd6716: data = 8'h80;
            20'd6717: data = 8'h80;
            20'd6718: data = 8'h80;
            20'd6719: data = 8'h80;
            20'd6720: data = 8'h80;
            20'd6721: data = 8'h80;
            20'd6722: data = 8'h80;
            20'd6723: data = 8'h80;
            20'd6724: data = 8'h80;
            20'd6725: data = 8'h80;
            20'd6726: data = 8'h80;
            20'd6727: data = 8'h80;
            20'd6728: data = 8'h80;
            20'd6729: data = 8'h80;
            20'd6730: data = 8'h80;
            20'd6731: data = 8'h80;
            20'd6732: data = 8'h80;
            20'd6733: data = 8'h80;
            20'd6734: data = 8'h80;
            20'd6735: data = 8'h80;
            20'd6736: data = 8'h80;
            20'd6737: data = 8'h80;
            20'd6738: data = 8'h80;
            20'd6739: data = 8'h80;
            20'd6740: data = 8'h80;
            20'd6741: data = 8'h80;
            20'd6742: data = 8'h80;
            20'd6743: data = 8'h80;
            20'd6744: data = 8'h80;
            20'd6745: data = 8'h80;
            20'd6746: data = 8'h80;
            20'd6747: data = 8'h80;
            20'd6748: data = 8'h80;
            20'd6749: data = 8'h80;
            20'd6750: data = 8'h80;
            20'd6751: data = 8'h80;
            20'd6752: data = 8'h80;
            20'd6753: data = 8'h80;
            20'd6754: data = 8'h80;
            20'd6755: data = 8'h80;
            20'd6756: data = 8'h80;
            20'd6757: data = 8'h80;
            20'd6758: data = 8'h80;
            20'd6759: data = 8'h80;
            20'd6760: data = 8'h80;
            20'd6761: data = 8'h80;
            20'd6762: data = 8'h80;
            20'd6763: data = 8'h80;
            20'd6764: data = 8'h80;
            20'd6765: data = 8'h80;
            20'd6766: data = 8'h80;
            20'd6767: data = 8'h80;
            20'd6768: data = 8'h80;
            20'd6769: data = 8'h80;
            20'd6770: data = 8'h80;
            20'd6771: data = 8'h80;
            20'd6772: data = 8'h80;
            20'd6773: data = 8'h80;
            20'd6774: data = 8'h80;
            20'd6775: data = 8'h80;
            20'd6776: data = 8'h80;
            20'd6777: data = 8'h80;
            20'd6778: data = 8'h80;
            20'd6779: data = 8'h80;
            20'd6780: data = 8'h80;
            20'd6781: data = 8'h80;
            20'd6782: data = 8'h80;
            20'd6783: data = 8'h80;
            20'd6784: data = 8'h80;
            20'd6785: data = 8'h80;
            20'd6786: data = 8'h80;
            20'd6787: data = 8'h80;
            20'd6788: data = 8'h80;
            20'd6789: data = 8'h80;
            20'd6790: data = 8'h80;
            20'd6791: data = 8'h80;
            20'd6792: data = 8'h80;
            20'd6793: data = 8'h80;
            20'd6794: data = 8'h80;
            20'd6795: data = 8'h80;
            20'd6796: data = 8'h80;
            20'd6797: data = 8'h80;
            20'd6798: data = 8'h80;
            20'd6799: data = 8'h80;
            20'd6800: data = 8'h80;
            20'd6801: data = 8'h80;
            20'd6802: data = 8'h80;
            20'd6803: data = 8'h80;
            20'd6804: data = 8'h80;
            20'd6805: data = 8'h80;
            20'd6806: data = 8'h80;
            20'd6807: data = 8'h80;
            20'd6808: data = 8'h80;
            20'd6809: data = 8'h80;
            20'd6810: data = 8'h80;
            20'd6811: data = 8'h80;
            20'd6812: data = 8'h80;
            20'd6813: data = 8'h80;
            20'd6814: data = 8'h80;
            20'd6815: data = 8'h80;
            20'd6816: data = 8'h80;
            20'd6817: data = 8'h80;
            20'd6818: data = 8'h80;
            20'd6819: data = 8'h80;
            20'd6820: data = 8'h80;
            20'd6821: data = 8'h80;
            20'd6822: data = 8'h80;
            20'd6823: data = 8'h80;
            20'd6824: data = 8'h80;
            20'd6825: data = 8'h80;
            20'd6826: data = 8'h80;
            20'd6827: data = 8'h80;
            20'd6828: data = 8'h80;
            20'd6829: data = 8'h80;
            20'd6830: data = 8'h80;
            20'd6831: data = 8'h80;
            20'd6832: data = 8'h80;
            20'd6833: data = 8'h80;
            20'd6834: data = 8'h80;
            20'd6835: data = 8'h80;
            20'd6836: data = 8'h80;
            20'd6837: data = 8'h80;
            20'd6838: data = 8'h80;
            20'd6839: data = 8'h80;
            20'd6840: data = 8'h80;
            20'd6841: data = 8'h80;
            20'd6842: data = 8'h80;
            20'd6843: data = 8'h80;
            20'd6844: data = 8'h80;
            20'd6845: data = 8'h80;
            20'd6846: data = 8'h80;
            20'd6847: data = 8'h80;
            20'd6848: data = 8'h80;
            20'd6849: data = 8'h80;
            20'd6850: data = 8'h80;
            20'd6851: data = 8'h80;
            20'd6852: data = 8'h80;
            20'd6853: data = 8'h80;
            20'd6854: data = 8'h80;
            20'd6855: data = 8'h80;
            20'd6856: data = 8'h80;
            20'd6857: data = 8'h80;
            20'd6858: data = 8'h80;
            20'd6859: data = 8'h80;
            20'd6860: data = 8'h80;
            20'd6861: data = 8'h80;
            20'd6862: data = 8'h80;
            20'd6863: data = 8'h80;
            20'd6864: data = 8'h80;
            20'd6865: data = 8'h80;
            20'd6866: data = 8'h80;
            20'd6867: data = 8'h80;
            20'd6868: data = 8'h80;
            20'd6869: data = 8'h80;
            20'd6870: data = 8'h80;
            20'd6871: data = 8'h80;
            20'd6872: data = 8'h80;
            20'd6873: data = 8'h80;
            20'd6874: data = 8'h80;
            20'd6875: data = 8'h80;
            20'd6876: data = 8'h80;
            20'd6877: data = 8'h80;
            20'd6878: data = 8'h80;
            20'd6879: data = 8'h80;
            20'd6880: data = 8'h80;
            20'd6881: data = 8'h80;
            20'd6882: data = 8'h80;
            20'd6883: data = 8'h80;
            20'd6884: data = 8'h80;
            20'd6885: data = 8'h80;
            20'd6886: data = 8'h80;
            20'd6887: data = 8'h80;
            20'd6888: data = 8'h80;
            20'd6889: data = 8'h80;
            20'd6890: data = 8'h80;
            20'd6891: data = 8'h80;
            20'd6892: data = 8'h80;
            20'd6893: data = 8'h80;
            20'd6894: data = 8'h80;
            20'd6895: data = 8'h80;
            20'd6896: data = 8'h80;
            20'd6897: data = 8'h80;
            20'd6898: data = 8'h80;
            20'd6899: data = 8'h80;
            20'd6900: data = 8'h80;
            20'd6901: data = 8'h80;
            20'd6902: data = 8'h80;
            20'd6903: data = 8'h80;
            20'd6904: data = 8'h80;
            20'd6905: data = 8'h80;
            20'd6906: data = 8'h80;
            20'd6907: data = 8'h80;
            20'd6908: data = 8'h80;
            20'd6909: data = 8'h80;
            20'd6910: data = 8'h80;
            20'd6911: data = 8'h80;
            20'd6912: data = 8'h80;
            20'd6913: data = 8'h80;
            20'd6914: data = 8'h80;
            20'd6915: data = 8'h80;
            20'd6916: data = 8'h80;
            20'd6917: data = 8'h80;
            20'd6918: data = 8'h80;
            20'd6919: data = 8'h80;
            20'd6920: data = 8'h80;
            20'd6921: data = 8'h80;
            20'd6922: data = 8'h80;
            20'd6923: data = 8'h80;
            20'd6924: data = 8'h80;
            20'd6925: data = 8'h80;
            20'd6926: data = 8'h80;
            20'd6927: data = 8'h80;
            20'd6928: data = 8'h80;
            20'd6929: data = 8'h80;
            20'd6930: data = 8'h80;
            20'd6931: data = 8'h80;
            20'd6932: data = 8'h80;
            20'd6933: data = 8'h80;
            20'd6934: data = 8'h80;
            20'd6935: data = 8'h80;
            20'd6936: data = 8'h80;
            20'd6937: data = 8'h80;
            20'd6938: data = 8'h80;
            20'd6939: data = 8'h80;
            20'd6940: data = 8'h80;
            20'd6941: data = 8'h80;
            20'd6942: data = 8'h80;
            20'd6943: data = 8'h80;
            20'd6944: data = 8'h80;
            20'd6945: data = 8'h80;
            20'd6946: data = 8'h80;
            20'd6947: data = 8'h80;
            20'd6948: data = 8'h80;
            20'd6949: data = 8'h80;
            20'd6950: data = 8'h80;
            20'd6951: data = 8'h80;
            20'd6952: data = 8'h80;
            20'd6953: data = 8'h80;
            20'd6954: data = 8'h80;
            20'd6955: data = 8'h80;
            20'd6956: data = 8'h80;
            20'd6957: data = 8'h80;
            20'd6958: data = 8'h80;
            20'd6959: data = 8'h80;
            20'd6960: data = 8'h80;
            20'd6961: data = 8'h80;
            20'd6962: data = 8'h80;
            20'd6963: data = 8'h80;
            20'd6964: data = 8'h80;
            20'd6965: data = 8'h80;
            20'd6966: data = 8'h80;
            20'd6967: data = 8'h80;
            20'd6968: data = 8'h80;
            20'd6969: data = 8'h80;
            20'd6970: data = 8'h80;
            20'd6971: data = 8'h80;
            20'd6972: data = 8'h80;
            20'd6973: data = 8'h80;
            20'd6974: data = 8'h80;
            20'd6975: data = 8'h80;
            20'd6976: data = 8'h80;
            20'd6977: data = 8'h80;
            20'd6978: data = 8'h80;
            20'd6979: data = 8'h80;
            20'd6980: data = 8'h80;
            20'd6981: data = 8'h80;
            20'd6982: data = 8'h80;
            20'd6983: data = 8'h80;
            20'd6984: data = 8'h80;
            20'd6985: data = 8'h80;
            20'd6986: data = 8'h80;
            20'd6987: data = 8'h80;
            20'd6988: data = 8'h80;
            20'd6989: data = 8'h80;
            20'd6990: data = 8'h80;
            20'd6991: data = 8'h80;
            20'd6992: data = 8'h80;
            20'd6993: data = 8'h80;
            20'd6994: data = 8'h80;
            20'd6995: data = 8'h80;
            20'd6996: data = 8'h80;
            20'd6997: data = 8'h80;
            20'd6998: data = 8'h80;
            20'd6999: data = 8'h80;
            20'd7000: data = 8'h80;
            20'd7001: data = 8'h80;
            20'd7002: data = 8'h80;
            20'd7003: data = 8'h80;
            20'd7004: data = 8'h80;
            20'd7005: data = 8'h80;
            20'd7006: data = 8'h80;
            20'd7007: data = 8'h80;
            20'd7008: data = 8'h80;
            20'd7009: data = 8'h80;
            20'd7010: data = 8'h80;
            20'd7011: data = 8'h80;
            20'd7012: data = 8'h80;
            20'd7013: data = 8'h80;
            20'd7014: data = 8'h80;
            20'd7015: data = 8'h80;
            20'd7016: data = 8'h80;
            20'd7017: data = 8'h80;
            20'd7018: data = 8'h80;
            20'd7019: data = 8'h80;
            20'd7020: data = 8'h80;
            20'd7021: data = 8'h80;
            20'd7022: data = 8'h80;
            20'd7023: data = 8'h80;
            20'd7024: data = 8'h80;
            20'd7025: data = 8'h80;
            20'd7026: data = 8'h80;
            20'd7027: data = 8'h80;
            20'd7028: data = 8'h80;
            20'd7029: data = 8'h80;
            20'd7030: data = 8'h80;
            20'd7031: data = 8'h80;
            20'd7032: data = 8'h80;
            20'd7033: data = 8'h80;
            20'd7034: data = 8'h80;
            20'd7035: data = 8'h80;
            20'd7036: data = 8'h80;
            20'd7037: data = 8'h80;
            20'd7038: data = 8'h80;
            20'd7039: data = 8'h80;
            20'd7040: data = 8'h80;
            20'd7041: data = 8'h80;
            20'd7042: data = 8'h80;
            20'd7043: data = 8'h80;
            20'd7044: data = 8'h80;
            20'd7045: data = 8'h80;
            20'd7046: data = 8'h80;
            20'd7047: data = 8'h80;
            20'd7048: data = 8'h80;
            20'd7049: data = 8'h80;
            20'd7050: data = 8'h80;
            20'd7051: data = 8'h80;
            20'd7052: data = 8'h80;
            20'd7053: data = 8'h80;
            20'd7054: data = 8'h80;
            20'd7055: data = 8'h80;
            20'd7056: data = 8'h80;
            20'd7057: data = 8'h80;
            20'd7058: data = 8'h80;
            20'd7059: data = 8'h80;
            20'd7060: data = 8'h80;
            20'd7061: data = 8'h80;
            20'd7062: data = 8'h80;
            20'd7063: data = 8'h80;
            20'd7064: data = 8'h80;
            20'd7065: data = 8'h80;
            20'd7066: data = 8'h80;
            20'd7067: data = 8'h80;
            20'd7068: data = 8'h80;
            20'd7069: data = 8'h80;
            20'd7070: data = 8'h80;
            20'd7071: data = 8'h80;
            20'd7072: data = 8'h80;
            20'd7073: data = 8'h80;
            20'd7074: data = 8'h80;
            20'd7075: data = 8'h80;
            20'd7076: data = 8'h80;
            20'd7077: data = 8'h80;
            20'd7078: data = 8'h80;
            20'd7079: data = 8'h80;
            20'd7080: data = 8'h80;
            20'd7081: data = 8'h80;
            20'd7082: data = 8'h80;
            20'd7083: data = 8'h80;
            20'd7084: data = 8'h80;
            20'd7085: data = 8'h80;
            20'd7086: data = 8'h80;
            20'd7087: data = 8'h80;
            20'd7088: data = 8'h80;
            20'd7089: data = 8'h80;
            20'd7090: data = 8'h80;
            20'd7091: data = 8'h80;
            20'd7092: data = 8'h80;
            20'd7093: data = 8'h80;
            20'd7094: data = 8'h80;
            20'd7095: data = 8'h80;
            20'd7096: data = 8'h80;
            20'd7097: data = 8'h80;
            20'd7098: data = 8'h80;
            20'd7099: data = 8'h80;
            20'd7100: data = 8'h80;
            20'd7101: data = 8'h80;
            20'd7102: data = 8'h80;
            20'd7103: data = 8'h80;
            20'd7104: data = 8'h80;
            20'd7105: data = 8'h80;
            20'd7106: data = 8'h80;
            20'd7107: data = 8'h80;
            20'd7108: data = 8'h80;
            20'd7109: data = 8'h80;
            20'd7110: data = 8'h80;
            20'd7111: data = 8'h80;
            20'd7112: data = 8'h80;
            20'd7113: data = 8'h80;
            20'd7114: data = 8'h80;
            20'd7115: data = 8'h80;
            20'd7116: data = 8'h80;
            20'd7117: data = 8'h80;
            20'd7118: data = 8'h80;
            20'd7119: data = 8'h80;
            20'd7120: data = 8'h80;
            20'd7121: data = 8'h80;
            20'd7122: data = 8'h80;
            20'd7123: data = 8'h80;
            20'd7124: data = 8'h80;
            20'd7125: data = 8'h80;
            20'd7126: data = 8'h80;
            20'd7127: data = 8'h80;
            20'd7128: data = 8'h80;
            20'd7129: data = 8'h80;
            20'd7130: data = 8'h80;
            20'd7131: data = 8'h80;
            20'd7132: data = 8'h80;
            20'd7133: data = 8'h80;
            20'd7134: data = 8'h80;
            20'd7135: data = 8'h80;
            20'd7136: data = 8'h80;
            20'd7137: data = 8'h80;
            20'd7138: data = 8'h80;
            20'd7139: data = 8'h80;
            20'd7140: data = 8'h80;
            20'd7141: data = 8'h80;
            20'd7142: data = 8'h80;
            20'd7143: data = 8'h80;
            20'd7144: data = 8'h80;
            20'd7145: data = 8'h80;
            20'd7146: data = 8'h80;
            20'd7147: data = 8'h80;
            20'd7148: data = 8'h80;
            20'd7149: data = 8'h80;
            20'd7150: data = 8'h80;
            20'd7151: data = 8'h80;
            20'd7152: data = 8'h80;
            20'd7153: data = 8'h80;
            20'd7154: data = 8'h80;
            20'd7155: data = 8'h80;
            20'd7156: data = 8'h80;
            20'd7157: data = 8'h80;
            20'd7158: data = 8'h80;
            20'd7159: data = 8'h80;
            20'd7160: data = 8'h80;
            20'd7161: data = 8'h80;
            20'd7162: data = 8'h80;
            20'd7163: data = 8'h80;
            20'd7164: data = 8'h80;
            20'd7165: data = 8'h80;
            20'd7166: data = 8'h80;
            20'd7167: data = 8'h80;
            20'd7168: data = 8'h80;
            20'd7169: data = 8'h80;
            20'd7170: data = 8'h80;
            20'd7171: data = 8'h80;
            20'd7172: data = 8'h80;
            20'd7173: data = 8'h80;
            20'd7174: data = 8'h80;
            20'd7175: data = 8'h80;
            20'd7176: data = 8'h80;
            20'd7177: data = 8'h80;
            20'd7178: data = 8'h80;
            20'd7179: data = 8'h80;
            20'd7180: data = 8'h80;
            20'd7181: data = 8'h80;
            20'd7182: data = 8'h80;
            20'd7183: data = 8'h80;
            20'd7184: data = 8'h80;
            20'd7185: data = 8'h80;
            20'd7186: data = 8'h80;
            20'd7187: data = 8'h80;
            20'd7188: data = 8'h80;
            20'd7189: data = 8'h80;
            20'd7190: data = 8'h80;
            20'd7191: data = 8'h80;
            20'd7192: data = 8'h80;
            20'd7193: data = 8'h80;
            20'd7194: data = 8'h80;
            20'd7195: data = 8'h80;
            20'd7196: data = 8'h80;
            20'd7197: data = 8'h80;
            20'd7198: data = 8'h80;
            20'd7199: data = 8'h80;
            20'd7200: data = 8'h80;
            20'd7201: data = 8'h80;
            20'd7202: data = 8'h80;
            20'd7203: data = 8'h80;
            20'd7204: data = 8'h80;
            20'd7205: data = 8'h80;
            20'd7206: data = 8'h80;
            20'd7207: data = 8'h80;
            20'd7208: data = 8'h80;
            20'd7209: data = 8'h80;
            20'd7210: data = 8'h80;
            20'd7211: data = 8'h80;
            20'd7212: data = 8'h80;
            20'd7213: data = 8'h80;
            20'd7214: data = 8'h80;
            20'd7215: data = 8'h80;
            20'd7216: data = 8'h80;
            20'd7217: data = 8'h80;
            20'd7218: data = 8'h80;
            20'd7219: data = 8'h80;
            20'd7220: data = 8'h80;
            20'd7221: data = 8'h80;
            20'd7222: data = 8'h80;
            20'd7223: data = 8'h80;
            20'd7224: data = 8'h80;
            20'd7225: data = 8'h80;
            20'd7226: data = 8'h80;
            20'd7227: data = 8'h80;
            20'd7228: data = 8'h80;
            20'd7229: data = 8'h80;
            20'd7230: data = 8'h80;
            20'd7231: data = 8'h80;
            20'd7232: data = 8'h80;
            20'd7233: data = 8'h80;
            20'd7234: data = 8'h80;
            20'd7235: data = 8'h80;
            20'd7236: data = 8'h80;
            20'd7237: data = 8'h80;
            20'd7238: data = 8'h80;
            20'd7239: data = 8'h80;
            20'd7240: data = 8'h80;
            20'd7241: data = 8'h80;
            20'd7242: data = 8'h80;
            20'd7243: data = 8'h80;
            20'd7244: data = 8'h80;
            20'd7245: data = 8'h80;
            20'd7246: data = 8'h80;
            20'd7247: data = 8'h80;
            20'd7248: data = 8'h80;
            20'd7249: data = 8'h80;
            20'd7250: data = 8'h80;
            20'd7251: data = 8'h80;
            20'd7252: data = 8'h80;
            20'd7253: data = 8'h80;
            20'd7254: data = 8'h80;
            20'd7255: data = 8'h80;
            20'd7256: data = 8'h80;
            20'd7257: data = 8'h80;
            20'd7258: data = 8'h80;
            20'd7259: data = 8'h80;
            20'd7260: data = 8'h80;
            20'd7261: data = 8'h80;
            20'd7262: data = 8'h80;
            20'd7263: data = 8'h80;
            20'd7264: data = 8'h80;
            20'd7265: data = 8'h80;
            20'd7266: data = 8'h80;
            20'd7267: data = 8'h80;
            20'd7268: data = 8'h80;
            20'd7269: data = 8'h80;
            20'd7270: data = 8'h80;
            20'd7271: data = 8'h80;
            20'd7272: data = 8'h80;
            20'd7273: data = 8'h80;
            20'd7274: data = 8'h80;
            20'd7275: data = 8'h80;
            20'd7276: data = 8'h80;
            20'd7277: data = 8'h80;
            20'd7278: data = 8'h80;
            20'd7279: data = 8'h80;
            20'd7280: data = 8'h80;
            20'd7281: data = 8'h80;
            20'd7282: data = 8'h80;
            20'd7283: data = 8'h80;
            20'd7284: data = 8'h80;
            20'd7285: data = 8'h80;
            20'd7286: data = 8'h80;
            20'd7287: data = 8'h80;
            20'd7288: data = 8'h80;
            20'd7289: data = 8'h80;
            20'd7290: data = 8'h80;
            20'd7291: data = 8'h80;
            20'd7292: data = 8'h80;
            20'd7293: data = 8'h80;
            20'd7294: data = 8'h80;
            20'd7295: data = 8'h80;
            20'd7296: data = 8'h80;
            20'd7297: data = 8'h80;
            20'd7298: data = 8'h80;
            20'd7299: data = 8'h80;
            20'd7300: data = 8'h80;
            20'd7301: data = 8'h80;
            20'd7302: data = 8'h80;
            20'd7303: data = 8'h80;
            20'd7304: data = 8'h80;
            20'd7305: data = 8'h80;
            20'd7306: data = 8'h80;
            20'd7307: data = 8'h80;
            20'd7308: data = 8'h80;
            20'd7309: data = 8'h80;
            20'd7310: data = 8'h80;
            20'd7311: data = 8'h80;
            20'd7312: data = 8'h80;
            20'd7313: data = 8'h80;
            20'd7314: data = 8'h80;
            20'd7315: data = 8'h80;
            20'd7316: data = 8'h80;
            20'd7317: data = 8'h80;
            20'd7318: data = 8'h80;
            20'd7319: data = 8'h80;
            20'd7320: data = 8'h80;
            20'd7321: data = 8'h80;
            20'd7322: data = 8'h80;
            20'd7323: data = 8'h80;
            20'd7324: data = 8'h80;
            20'd7325: data = 8'h80;
            20'd7326: data = 8'h80;
            20'd7327: data = 8'h80;
            20'd7328: data = 8'h80;
            20'd7329: data = 8'h80;
            20'd7330: data = 8'h80;
            20'd7331: data = 8'h80;
            20'd7332: data = 8'h80;
            20'd7333: data = 8'h80;
            20'd7334: data = 8'h80;
            20'd7335: data = 8'h80;
            20'd7336: data = 8'h80;
            20'd7337: data = 8'h80;
            20'd7338: data = 8'h80;
            20'd7339: data = 8'h80;
            20'd7340: data = 8'h80;
            20'd7341: data = 8'h80;
            20'd7342: data = 8'h80;
            20'd7343: data = 8'h80;
            20'd7344: data = 8'h80;
            20'd7345: data = 8'h80;
            20'd7346: data = 8'h80;
            20'd7347: data = 8'h80;
            20'd7348: data = 8'h80;
            20'd7349: data = 8'h80;
            20'd7350: data = 8'h80;
            20'd7351: data = 8'h80;
            20'd7352: data = 8'h80;
            20'd7353: data = 8'h80;
            20'd7354: data = 8'h80;
            20'd7355: data = 8'h80;
            20'd7356: data = 8'h80;
            20'd7357: data = 8'h80;
            20'd7358: data = 8'h80;
            20'd7359: data = 8'h80;
            20'd7360: data = 8'h80;
            20'd7361: data = 8'h80;
            20'd7362: data = 8'h80;
            20'd7363: data = 8'h80;
            20'd7364: data = 8'h80;
            20'd7365: data = 8'h80;
            20'd7366: data = 8'h80;
            20'd7367: data = 8'h80;
            20'd7368: data = 8'h80;
            20'd7369: data = 8'h80;
            20'd7370: data = 8'h80;
            20'd7371: data = 8'h80;
            20'd7372: data = 8'h80;
            20'd7373: data = 8'h80;
            20'd7374: data = 8'h80;
            20'd7375: data = 8'h80;
            20'd7376: data = 8'h80;
            20'd7377: data = 8'h80;
            20'd7378: data = 8'h80;
            20'd7379: data = 8'h80;
            20'd7380: data = 8'h80;
            20'd7381: data = 8'h80;
            20'd7382: data = 8'h80;
            20'd7383: data = 8'h80;
            20'd7384: data = 8'h80;
            20'd7385: data = 8'h80;
            20'd7386: data = 8'h80;
            20'd7387: data = 8'h80;
            20'd7388: data = 8'h80;
            20'd7389: data = 8'h80;
            20'd7390: data = 8'h80;
            20'd7391: data = 8'h80;
            20'd7392: data = 8'h80;
            20'd7393: data = 8'h80;
            20'd7394: data = 8'h80;
            20'd7395: data = 8'h80;
            20'd7396: data = 8'h80;
            20'd7397: data = 8'h80;
            20'd7398: data = 8'h80;
            20'd7399: data = 8'h80;
            20'd7400: data = 8'h80;
            20'd7401: data = 8'h80;
            20'd7402: data = 8'h80;
            20'd7403: data = 8'h80;
            20'd7404: data = 8'h80;
            20'd7405: data = 8'h80;
            20'd7406: data = 8'h80;
            20'd7407: data = 8'h80;
            20'd7408: data = 8'h80;
            20'd7409: data = 8'h80;
            20'd7410: data = 8'h80;
            20'd7411: data = 8'h80;
            20'd7412: data = 8'h80;
            20'd7413: data = 8'h80;
            20'd7414: data = 8'h80;
            20'd7415: data = 8'h80;
            20'd7416: data = 8'h80;
            20'd7417: data = 8'h80;
            20'd7418: data = 8'h80;
            20'd7419: data = 8'h80;
            20'd7420: data = 8'h80;
            20'd7421: data = 8'h80;
            20'd7422: data = 8'h80;
            20'd7423: data = 8'h80;
            20'd7424: data = 8'h80;
            20'd7425: data = 8'h80;
            20'd7426: data = 8'h80;
            20'd7427: data = 8'h80;
            20'd7428: data = 8'h80;
            20'd7429: data = 8'h80;
            20'd7430: data = 8'h80;
            20'd7431: data = 8'h80;
            20'd7432: data = 8'h80;
            20'd7433: data = 8'h80;
            20'd7434: data = 8'h80;
            20'd7435: data = 8'h80;
            20'd7436: data = 8'h80;
            20'd7437: data = 8'h80;
            20'd7438: data = 8'h80;
            20'd7439: data = 8'h80;
            20'd7440: data = 8'h80;
            20'd7441: data = 8'h80;
            20'd7442: data = 8'h80;
            20'd7443: data = 8'h80;
            20'd7444: data = 8'h80;
            20'd7445: data = 8'h80;
            20'd7446: data = 8'h80;
            20'd7447: data = 8'h80;
            20'd7448: data = 8'h80;
            20'd7449: data = 8'h80;
            20'd7450: data = 8'h80;
            20'd7451: data = 8'h80;
            20'd7452: data = 8'h80;
            20'd7453: data = 8'h80;
            20'd7454: data = 8'h80;
            20'd7455: data = 8'h80;
            20'd7456: data = 8'h80;
            20'd7457: data = 8'h80;
            20'd7458: data = 8'h80;
            20'd7459: data = 8'h80;
            20'd7460: data = 8'h80;
            20'd7461: data = 8'h80;
            20'd7462: data = 8'h80;
            20'd7463: data = 8'h80;
            20'd7464: data = 8'h80;
            20'd7465: data = 8'h80;
            20'd7466: data = 8'h80;
            20'd7467: data = 8'h80;
            20'd7468: data = 8'h80;
            20'd7469: data = 8'h80;
            20'd7470: data = 8'h80;
            20'd7471: data = 8'h80;
            20'd7472: data = 8'h80;
            20'd7473: data = 8'h80;
            20'd7474: data = 8'h80;
            20'd7475: data = 8'h80;
            20'd7476: data = 8'h80;
            20'd7477: data = 8'h80;
            20'd7478: data = 8'h80;
            20'd7479: data = 8'h80;
            20'd7480: data = 8'h80;
            20'd7481: data = 8'h80;
            20'd7482: data = 8'h80;
            20'd7483: data = 8'h80;
            20'd7484: data = 8'h80;
            20'd7485: data = 8'h80;
            20'd7486: data = 8'h80;
            20'd7487: data = 8'h80;
            20'd7488: data = 8'h80;
            20'd7489: data = 8'h80;
            20'd7490: data = 8'h80;
            20'd7491: data = 8'h80;
            20'd7492: data = 8'h80;
            20'd7493: data = 8'h80;
            20'd7494: data = 8'h80;
            20'd7495: data = 8'h80;
            20'd7496: data = 8'h80;
            20'd7497: data = 8'h80;
            20'd7498: data = 8'h80;
            20'd7499: data = 8'h80;
            20'd7500: data = 8'h80;
            20'd7501: data = 8'h80;
            20'd7502: data = 8'h80;
            20'd7503: data = 8'h80;
            20'd7504: data = 8'h80;
            20'd7505: data = 8'h80;
            20'd7506: data = 8'h80;
            20'd7507: data = 8'h80;
            20'd7508: data = 8'h80;
            20'd7509: data = 8'h80;
            20'd7510: data = 8'h80;
            20'd7511: data = 8'h80;
            20'd7512: data = 8'h80;
            20'd7513: data = 8'h80;
            20'd7514: data = 8'h80;
            20'd7515: data = 8'h80;
            20'd7516: data = 8'h80;
            20'd7517: data = 8'h80;
            20'd7518: data = 8'h80;
            20'd7519: data = 8'h80;
            20'd7520: data = 8'h80;
            20'd7521: data = 8'h80;
            20'd7522: data = 8'h80;
            20'd7523: data = 8'h80;
            20'd7524: data = 8'h80;
            20'd7525: data = 8'h80;
            20'd7526: data = 8'h80;
            20'd7527: data = 8'h80;
            20'd7528: data = 8'h80;
            20'd7529: data = 8'h80;
            20'd7530: data = 8'h80;
            20'd7531: data = 8'h80;
            20'd7532: data = 8'h80;
            20'd7533: data = 8'h80;
            20'd7534: data = 8'h80;
            20'd7535: data = 8'h80;
            20'd7536: data = 8'h80;
            20'd7537: data = 8'h80;
            20'd7538: data = 8'h80;
            20'd7539: data = 8'h80;
            20'd7540: data = 8'h80;
            20'd7541: data = 8'h80;
            20'd7542: data = 8'h80;
            20'd7543: data = 8'h80;
            20'd7544: data = 8'h80;
            20'd7545: data = 8'h80;
            20'd7546: data = 8'h80;
            20'd7547: data = 8'h80;
            20'd7548: data = 8'h80;
            20'd7549: data = 8'h80;
            20'd7550: data = 8'h80;
            20'd7551: data = 8'h80;
            20'd7552: data = 8'h80;
            20'd7553: data = 8'h80;
            20'd7554: data = 8'h80;
            20'd7555: data = 8'h80;
            20'd7556: data = 8'h80;
            20'd7557: data = 8'h80;
            20'd7558: data = 8'h80;
            20'd7559: data = 8'h80;
            20'd7560: data = 8'h80;
            20'd7561: data = 8'h80;
            20'd7562: data = 8'h80;
            20'd7563: data = 8'h80;
            20'd7564: data = 8'h80;
            20'd7565: data = 8'h80;
            20'd7566: data = 8'h80;
            20'd7567: data = 8'h80;
            20'd7568: data = 8'h80;
            20'd7569: data = 8'h80;
            20'd7570: data = 8'h80;
            20'd7571: data = 8'h80;
            20'd7572: data = 8'h80;
            20'd7573: data = 8'h80;
            20'd7574: data = 8'h80;
            20'd7575: data = 8'h80;
            20'd7576: data = 8'h80;
            20'd7577: data = 8'h80;
            20'd7578: data = 8'h80;
            20'd7579: data = 8'h80;
            20'd7580: data = 8'h80;
            20'd7581: data = 8'h80;
            20'd7582: data = 8'h80;
            20'd7583: data = 8'h80;
            20'd7584: data = 8'h80;
            20'd7585: data = 8'h80;
            20'd7586: data = 8'h80;
            20'd7587: data = 8'h80;
            20'd7588: data = 8'h80;
            20'd7589: data = 8'h80;
            20'd7590: data = 8'h80;
            20'd7591: data = 8'h80;
            20'd7592: data = 8'h80;
            20'd7593: data = 8'h80;
            20'd7594: data = 8'h80;
            20'd7595: data = 8'h80;
            20'd7596: data = 8'h80;
            20'd7597: data = 8'h80;
            20'd7598: data = 8'h80;
            20'd7599: data = 8'h80;
            20'd7600: data = 8'h80;
            20'd7601: data = 8'h80;
            20'd7602: data = 8'h80;
            20'd7603: data = 8'h80;
            20'd7604: data = 8'h80;
            20'd7605: data = 8'h80;
            20'd7606: data = 8'h80;
            20'd7607: data = 8'h80;
            20'd7608: data = 8'h80;
            20'd7609: data = 8'h80;
            20'd7610: data = 8'h80;
            20'd7611: data = 8'h80;
            20'd7612: data = 8'h80;
            20'd7613: data = 8'h80;
            20'd7614: data = 8'h80;
            20'd7615: data = 8'h80;
            20'd7616: data = 8'h80;
            20'd7617: data = 8'h80;
            20'd7618: data = 8'h80;
            20'd7619: data = 8'h80;
            20'd7620: data = 8'h80;
            20'd7621: data = 8'h80;
            20'd7622: data = 8'h80;
            20'd7623: data = 8'h80;
            20'd7624: data = 8'h80;
            20'd7625: data = 8'h80;
            20'd7626: data = 8'h80;
            20'd7627: data = 8'h80;
            20'd7628: data = 8'h80;
            20'd7629: data = 8'h80;
            20'd7630: data = 8'h80;
            20'd7631: data = 8'h80;
            20'd7632: data = 8'h80;
            20'd7633: data = 8'h80;
            20'd7634: data = 8'h80;
            20'd7635: data = 8'h80;
            20'd7636: data = 8'h80;
            20'd7637: data = 8'h80;
            20'd7638: data = 8'h80;
            20'd7639: data = 8'h80;
            20'd7640: data = 8'h80;
            20'd7641: data = 8'h80;
            20'd7642: data = 8'h80;
            20'd7643: data = 8'h80;
            20'd7644: data = 8'h80;
            20'd7645: data = 8'h80;
            20'd7646: data = 8'h80;
            20'd7647: data = 8'h80;
            20'd7648: data = 8'h80;
            20'd7649: data = 8'h80;
            20'd7650: data = 8'h80;
            20'd7651: data = 8'h80;
            20'd7652: data = 8'h80;
            20'd7653: data = 8'h80;
            20'd7654: data = 8'h80;
            20'd7655: data = 8'h80;
            20'd7656: data = 8'h80;
            20'd7657: data = 8'h80;
            20'd7658: data = 8'h80;
            20'd7659: data = 8'h80;
            20'd7660: data = 8'h80;
            20'd7661: data = 8'h80;
            20'd7662: data = 8'h80;
            20'd7663: data = 8'h80;
            20'd7664: data = 8'h80;
            20'd7665: data = 8'h80;
            20'd7666: data = 8'h80;
            20'd7667: data = 8'h80;
            20'd7668: data = 8'h80;
            20'd7669: data = 8'h80;
            20'd7670: data = 8'h80;
            20'd7671: data = 8'h80;
            20'd7672: data = 8'h80;
            20'd7673: data = 8'h80;
            20'd7674: data = 8'h80;
            20'd7675: data = 8'h80;
            20'd7676: data = 8'h80;
            20'd7677: data = 8'h80;
            20'd7678: data = 8'h80;
            20'd7679: data = 8'h80;
            20'd7680: data = 8'h80;
            20'd7681: data = 8'h80;
            20'd7682: data = 8'h80;
            20'd7683: data = 8'h80;
            20'd7684: data = 8'h80;
            20'd7685: data = 8'h80;
            20'd7686: data = 8'h80;
            20'd7687: data = 8'h80;
            20'd7688: data = 8'h80;
            20'd7689: data = 8'h80;
            20'd7690: data = 8'h80;
            20'd7691: data = 8'h80;
            20'd7692: data = 8'h80;
            20'd7693: data = 8'h80;
            20'd7694: data = 8'h80;
            20'd7695: data = 8'h80;
            20'd7696: data = 8'h80;
            20'd7697: data = 8'h80;
            20'd7698: data = 8'h80;
            20'd7699: data = 8'h80;
            20'd7700: data = 8'h80;
            20'd7701: data = 8'h80;
            20'd7702: data = 8'h80;
            20'd7703: data = 8'h80;
            20'd7704: data = 8'h80;
            20'd7705: data = 8'h80;
            20'd7706: data = 8'h80;
            20'd7707: data = 8'h80;
            20'd7708: data = 8'h80;
            20'd7709: data = 8'h80;
            20'd7710: data = 8'h80;
            20'd7711: data = 8'h80;
            20'd7712: data = 8'h80;
            20'd7713: data = 8'h80;
            20'd7714: data = 8'h80;
            20'd7715: data = 8'h80;
            20'd7716: data = 8'h80;
            20'd7717: data = 8'h80;
            20'd7718: data = 8'h80;
            20'd7719: data = 8'h80;
            20'd7720: data = 8'h80;
            20'd7721: data = 8'h80;
            20'd7722: data = 8'h80;
            20'd7723: data = 8'h80;
            20'd7724: data = 8'h80;
            20'd7725: data = 8'h80;
            20'd7726: data = 8'h80;
            20'd7727: data = 8'h80;
            20'd7728: data = 8'h80;
            20'd7729: data = 8'h80;
            20'd7730: data = 8'h80;
            20'd7731: data = 8'h80;
            20'd7732: data = 8'h80;
            20'd7733: data = 8'h80;
            20'd7734: data = 8'h80;
            20'd7735: data = 8'h80;
            20'd7736: data = 8'h80;
            20'd7737: data = 8'h80;
            20'd7738: data = 8'h80;
            20'd7739: data = 8'h80;
            20'd7740: data = 8'h80;
            20'd7741: data = 8'h80;
            20'd7742: data = 8'h80;
            20'd7743: data = 8'h80;
            20'd7744: data = 8'h80;
            20'd7745: data = 8'h80;
            20'd7746: data = 8'h80;
            20'd7747: data = 8'h80;
            20'd7748: data = 8'h80;
            20'd7749: data = 8'h80;
            20'd7750: data = 8'h80;
            20'd7751: data = 8'h80;
            20'd7752: data = 8'h80;
            20'd7753: data = 8'h80;
            20'd7754: data = 8'h80;
            20'd7755: data = 8'h80;
            20'd7756: data = 8'h80;
            20'd7757: data = 8'h80;
            20'd7758: data = 8'h80;
            20'd7759: data = 8'h80;
            20'd7760: data = 8'h80;
            20'd7761: data = 8'h80;
            20'd7762: data = 8'h80;
            20'd7763: data = 8'h80;
            20'd7764: data = 8'h80;
            20'd7765: data = 8'h80;
            20'd7766: data = 8'h80;
            20'd7767: data = 8'h80;
            20'd7768: data = 8'h80;
            20'd7769: data = 8'h80;
            20'd7770: data = 8'h80;
            20'd7771: data = 8'h80;
            20'd7772: data = 8'h80;
            20'd7773: data = 8'h80;
            20'd7774: data = 8'h80;
            20'd7775: data = 8'h80;
            20'd7776: data = 8'h80;
            20'd7777: data = 8'h80;
            20'd7778: data = 8'h80;
            20'd7779: data = 8'h80;
            20'd7780: data = 8'h80;
            20'd7781: data = 8'h80;
            20'd7782: data = 8'h80;
            20'd7783: data = 8'h80;
            20'd7784: data = 8'h80;
            20'd7785: data = 8'h80;
            20'd7786: data = 8'h80;
            20'd7787: data = 8'h80;
            20'd7788: data = 8'h80;
            20'd7789: data = 8'h80;
            20'd7790: data = 8'h80;
            20'd7791: data = 8'h80;
            20'd7792: data = 8'h80;
            20'd7793: data = 8'h80;
            20'd7794: data = 8'h80;
            20'd7795: data = 8'h80;
            20'd7796: data = 8'h80;
            20'd7797: data = 8'h80;
            20'd7798: data = 8'h80;
            20'd7799: data = 8'h80;
            20'd7800: data = 8'h80;
            20'd7801: data = 8'h80;
            20'd7802: data = 8'h80;
            20'd7803: data = 8'h80;
            20'd7804: data = 8'h80;
            20'd7805: data = 8'h80;
            20'd7806: data = 8'h80;
            20'd7807: data = 8'h80;
            20'd7808: data = 8'h80;
            20'd7809: data = 8'h80;
            20'd7810: data = 8'h80;
            20'd7811: data = 8'h80;
            20'd7812: data = 8'h80;
            20'd7813: data = 8'h80;
            20'd7814: data = 8'h80;
            20'd7815: data = 8'h80;
            20'd7816: data = 8'h80;
            20'd7817: data = 8'h80;
            20'd7818: data = 8'h80;
            20'd7819: data = 8'h80;
            20'd7820: data = 8'h80;
            20'd7821: data = 8'h80;
            20'd7822: data = 8'h80;
            20'd7823: data = 8'h80;
            20'd7824: data = 8'h80;
            20'd7825: data = 8'h80;
            20'd7826: data = 8'h80;
            20'd7827: data = 8'h80;
            20'd7828: data = 8'h80;
            20'd7829: data = 8'h80;
            20'd7830: data = 8'h80;
            20'd7831: data = 8'h80;
            20'd7832: data = 8'h80;
            20'd7833: data = 8'h80;
            20'd7834: data = 8'h80;
            20'd7835: data = 8'h80;
            20'd7836: data = 8'h80;
            20'd7837: data = 8'h80;
            20'd7838: data = 8'h80;
            20'd7839: data = 8'h80;
            20'd7840: data = 8'h80;
            20'd7841: data = 8'h80;
            20'd7842: data = 8'h80;
            20'd7843: data = 8'h80;
            20'd7844: data = 8'h80;
            20'd7845: data = 8'h80;
            20'd7846: data = 8'h80;
            20'd7847: data = 8'h80;
            20'd7848: data = 8'h80;
            20'd7849: data = 8'h80;
            20'd7850: data = 8'h80;
            20'd7851: data = 8'h80;
            20'd7852: data = 8'h80;
            20'd7853: data = 8'h80;
            20'd7854: data = 8'h80;
            20'd7855: data = 8'h80;
            20'd7856: data = 8'h80;
            20'd7857: data = 8'h80;
            20'd7858: data = 8'h80;
            20'd7859: data = 8'h80;
            20'd7860: data = 8'h80;
            20'd7861: data = 8'h80;
            20'd7862: data = 8'h80;
            20'd7863: data = 8'h80;
            20'd7864: data = 8'h80;
            20'd7865: data = 8'h80;
            20'd7866: data = 8'h80;
            20'd7867: data = 8'h80;
            20'd7868: data = 8'h80;
            20'd7869: data = 8'h80;
            20'd7870: data = 8'h80;
            20'd7871: data = 8'h80;
            20'd7872: data = 8'h80;
            20'd7873: data = 8'h80;
            20'd7874: data = 8'h80;
            20'd7875: data = 8'h80;
            20'd7876: data = 8'h80;
            20'd7877: data = 8'h80;
            20'd7878: data = 8'h80;
            20'd7879: data = 8'h80;
            20'd7880: data = 8'h80;
            20'd7881: data = 8'h80;
            20'd7882: data = 8'h80;
            20'd7883: data = 8'h80;
            20'd7884: data = 8'h80;
            20'd7885: data = 8'h80;
            20'd7886: data = 8'h80;
            20'd7887: data = 8'h80;
            20'd7888: data = 8'h80;
            20'd7889: data = 8'h80;
            20'd7890: data = 8'h80;
            20'd7891: data = 8'h80;
            20'd7892: data = 8'h80;
            20'd7893: data = 8'h80;
            20'd7894: data = 8'h80;
            20'd7895: data = 8'h80;
            20'd7896: data = 8'h80;
            20'd7897: data = 8'h80;
            20'd7898: data = 8'h80;
            20'd7899: data = 8'h80;
            20'd7900: data = 8'h80;
            20'd7901: data = 8'h80;
            20'd7902: data = 8'h80;
            20'd7903: data = 8'h80;
            20'd7904: data = 8'h80;
            20'd7905: data = 8'h80;
            20'd7906: data = 8'h80;
            20'd7907: data = 8'h80;
            20'd7908: data = 8'h80;
            20'd7909: data = 8'h80;
            20'd7910: data = 8'h80;
            20'd7911: data = 8'h80;
            20'd7912: data = 8'h80;
            20'd7913: data = 8'h80;
            20'd7914: data = 8'h80;
            20'd7915: data = 8'h80;
            20'd7916: data = 8'h80;
            20'd7917: data = 8'h80;
            20'd7918: data = 8'h80;
            20'd7919: data = 8'h80;
            20'd7920: data = 8'h80;
            20'd7921: data = 8'h80;
            20'd7922: data = 8'h80;
            20'd7923: data = 8'h80;
            20'd7924: data = 8'h80;
            20'd7925: data = 8'h80;
            20'd7926: data = 8'h80;
            20'd7927: data = 8'h80;
            20'd7928: data = 8'h80;
            20'd7929: data = 8'h80;
            20'd7930: data = 8'h80;
            20'd7931: data = 8'h80;
            20'd7932: data = 8'h80;
            20'd7933: data = 8'h80;
            20'd7934: data = 8'h80;
            20'd7935: data = 8'h80;
            20'd7936: data = 8'h80;
            20'd7937: data = 8'h80;
            default: data = 8'h00;
        endcase
    end
endmodule
